//TA demo pattern

`ifdef RTL
    `define CYCLE_TIME 20.0
`endif
`ifdef GATE
    `define CYCLE_TIME 20.0
`endif
`ifdef POST
    `define CYCLE_TIME 20.0
`endif
module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_weight, 
	out_mode,
    // Input signals
    out_valid, 
	out_code
);


`protected
_+/0I=I6[^QPeP=HeYag1)dI#I1K#4YGEH:IDUEQ._7#BWX;U;&W3)PQaPBKXOBG
b/]A;Y522,F-2P>4LN:78abWEQ)HPHM^CH+^aDDa6D>b@;US]JQf7fS0cY1UD8H-
/S4J\TI&3MVKX?ZSXgYSeTXM]>91dZeWLNM\dK@+\8;Zg?bSS)gdB&,^VYX7HZ#C
4N682]:L.JZD_1R8(RPSe?XM5$
`endprotected
output reg clk, rst_n, in_valid, out_mode;
output reg [2:0] in_weight;

input out_valid, out_code;


`protected
X>?5]I8-X&^S@R;1T;2N/L-#.9NaUMVJU6?dBXf>-79U-B5,#;(S6)L9-g_DXLBH
5_(c.6I&:-H/(A87?1&dOA._MK@,eJI&END?@(\HS7A12B=D?3/1=&Nc,^8P,8&:
7=OV0&HU_P\6A5I]#415DaD6a+LAN?U&VVZ&@gF.J+:5B6JC1JcWY;<fB0@-^5eW
:aR=H4g>&0HTH[3&GV0AYH.)17Q5=W8gb35DREO/;DT:eHc:F#aS>WVYEU>0#eP2
NYK:=GaGbLS1CU82cA(@La7:)[P?X:#@=QI9<XB;Dgc(1Z.&)52C)GAGP[:0JH@U
P[1AWJ92T(S;\0e,[bNZJV?Rd4-WOH.E.DRgGQM>g[.>#e4#Y,1J3\7HVEQ1NO)K
1S_@]G^-<N4[NK_45M;JOSA]2I_#P5fQD0,)V]BJ+-(dW)LQ[CeRA@1AON&QcbY<
e@8K#-7Y[KHcJ5NB)=;IVEgE;?a/_6If,UMX8HZT\dH3_H)VN8J3/&MgY_Q:1\;d
RK2VHYfF0TX=UAbG=D<?[Y407^63d<7VO=#,HPH/J3:O/-?N_YQIcZ,E3>bIbI\]
[d9^ceb2(28.2=62F_/dPJH<JMR9VE5eKVY4G=bNS@R]C@SeQB>4R<?X\-RbD-3Y
Zc4)<P^6=f8VP:Y=b\3V4;Z2ad6?YDcdc<>2g1P8+7a.=XXbA+GX\[AJ[3;6]MVc
]3R(XYf^cIY^)6ENMfZ=JMKE:L6f1QUI6Z@A/+=QR/3?Gg4+KV]bX&GaF7/5Ub&Q
g2H4JQ+-K_>U6T:Ng;##1)25IZHdEKJ<2OMIb5-<#D2)9\G+2EF8:^6NcBQS/BI-
ZW^K>QR8+]:^Q5JQ[M;SB9J:TR7_K\20M-6:dU)J4A@WJPZ1,?_[HG&d<>+7a3;:
#?FM4+G&)ffb]B_SW;R@8;Xe:3b:4;.#f@Yc,LGGHP(:/H?KeOCcMG<S-YO@Pe9Y
dEbe-UV5-a+a7VS4OBS>,-UV0A@3GIE\1YA0Eb?fOM=f+\B61^]\f6QefG>.]aNB
4dJR41B?aXRD[8G<AU?;-EKTAO>A60aa_YW#.\W>G:8;S+FS1-G.0T6AbK+Rf-35
6.G90OHBAA\Fg)4](E8=@EZd\@I2AY72g[UAGF2/?A#O/72^BfHRZb8=A3I4MI[3
6.5MeYe\9Z0:4V#;(O(Mac?O=UO3&ZMYV?].:[,5:E)7POcRAVE=ga\Ea_=._EON
J\d6O?&BKSK.,cV)AMP4(QSb[>-;4X:+f9/]0X1T5FX^QEaS:3^+<UfEJUN&@TDQ
L@_ZM>,)<b:JVMM>B?#DbK++]aA[;4fBG7.N;Y,;^3ML^Z=3;F/MPc,\8MU\cVJ1
RY@F.9e>.NP@0VJ5.>Tb^AfGU>D5/@Xc.c@&1^W^90ZMFWB6.9Q;+F1_a@RS.XbW
_AL_#KCQYL(/QaWcESD+[EGdOU^+]H;Q_TOLDbIU>LT;93\Ga1(/D/&.<e_<e)N9
I)fRL)#GR;E;eI[,Tg/bB2e6F+3>Cg0JVDL64^N./WU,M\/d7+;4W4e/Q&-W/RLL
7/S9WbHgIVB?DdM&R+c\N9NSGNBQ;31JIfXDY5?gV\YG2O1#dL,IM;W)NJ<dZ//c
R?>J=8g)^7B\7S.4-Da.R72N0H)5.fHIH4b<X]3#NKcb;8df+gfU:8ILUM6@2?#-
9\4GgV55;H&7EG7[eZfLHacQLc/=9D+eUH3B:ZYH:Y4+2PL@\QHK+6]WZA8e3#S)
P:ec5&;dg#XWA5Y_743dP9Y@&7+9a3M:)YC)S,57HTT@>WO_Q7S/DC?73bWU]OWL
<7f-HI?,/3^[//_0dGa#6(@7U7JUgRS#SDJLdA(V@^2<4gD;dCg8GPC3YebVMT1\
7NCEX2&/bP@3>SM@8OL7_0:V&&(NX(\(G1R&-+7:QQNNaE(KPF67MYa]KKMLN:_d
_:gQBQUKONb8>OK;?J(_\f@7b1ZeS/?,])75GT<b8[cY<N)6H=Bc7g>P=^J026<T
D4GM\TJ4V:0bJ-Ud-]Cg)T1b]dH>_R=4_bg;.fI^DQX86(62HXG+#f@0JM8NDMIE
CgY^H&8A(5>;QWXEFO9^e0T5BK&/[/C(L9MZL&A1UcV/4O=@WUS^cVJ5X/4^LERg
.c/2UcG<1./J2M7fHHM\L9f/))V:V.GfUN5DL0cKPgU]a;d?)+GgGI#=RDD55OF3
E<]=b<5FcR+2U]#gTJbZ&AI5BLab)bVP3S4O8?LWMXB6VD2QP4c)[:9@(7AF6I38
:SJF/dZ7:@&]+g9O^.b/RSO-EG-S[A.CVQ)KA#QI\0e<@7<865GGK]:G/365QQK>
CA^MN/W^X8;UE7)>9;<:7MP21K=L:P5]CL,S)b,&Z7g;BcaI50>MJc;4ID&2V@eW
Y^?:d_E,@2TQO?V8O^g9U/1RJK8C50OEL@dg)TX[C;??e;^a2Yc&P#:(8?8Ca++X
&d35Z-F#CO[_gcH_NS\[;;7QVO?I7:VKHNfXRJ&_166C8SPOU#Ff1;KSA.E<bND.
bMP,RYc6LO-H>ORS9R@)1S895c[YY^14:@Ka.PcD@X\.JdY-_PY@8[(4(Q<__=^C
S.I.TS(P^Q,XBH:d@E\df/3&.TN9JFeJ?ZeQWc7=W3:F;fO.E(E8YE\g38a+450.
10TP<-;8K87LXScC-3:aE((@=3PJ@8@#NLS^-.D9HRV8+>aXa1U_]>Q3NVD.B-XA
E:OaK3Q48GCQbRMN51XgeQK(9,\<^/Q2B?@5KW.U8]Ua6N6,3N-2HZ/-8)AQDTSH
@^/e0S7.0\Gfe1FOg=X56P1HE#6Q.RFO0Q1-=^_>J_M-aHfOZ39:B7W)G6@G1WSC
eHd@>3d=_fMGFP&QWO0Dbg5NSKQ0=/=YbFC6#QdQbM.G;^V,\^VIBL\6U@(QA65@
1Cgg@697Jff2]70L&Be/b_6=]0E3]dYd_]cWH<0.1Y;]61GO;86Q+D;]DdN]18X&
O/BWa@?QS@He11LQ1/S[NX-FA7df]X#\Hb>U42JL&CA_^NVgDGEYS8=;g[J\gYC3
G1PWe/)gHPMX><Ve,FVM)1cfQ7OBW]gB:>c;BT2\dcVN6I_A+f]WEC<(P0OEbJ.3
]NG+M@,(6.]Mb87BL+U(68Y>28GBX2-X<6G^=M=_fR+BZfga12F6ND2;ET@QQ2[M
=829[bI(9B;XQ-HKI4]M3WD^(89dI19?9cY&c[]ga1-PD9La#bC#dc\<.JT@2]-_
B&[T-cE]H,2PAIA&?+2&\)J,-WCSO0X]gIE]O;W5cB=_Ff1Ca>6SAe^e_N45FDU-
8BE9#FA[1C;TO+,V<;P9#=C(]PG[]P5@3GK><<2>;/ag@VVVe[4FMW1,TOUA?H6A
:4B]MR-DI9W+(;IY(W5PP?Rd&F7/7R>/eP3+bXEBDN59e-S]U4f3\3-+gf_>2(7]
L+P#b.]]=e&=&g[_g]=V#16(#DQTPa5C>XS?/0N8[B@0640J)MgP61bgdSXOW?Q#
Z);5d_&&Be\D&RKfS6OgLD-&XM7<-^;M&57-^H]R&c&[,9X^I<FUBeT&?=OCMVTf
.YJf78_;RdeFR1Dd[8:EU-OWfMXVdRL.?VHMP.=;4OKI=bbR1-_3)fP)1cK;3:Sc
67[;&]J>ZfBYc#]cA;KAYH8A]JCD+WXAeUH_af(fa#LG@A0\\?P,P67I#^KZ)faW
W>SP3\=Bg2(K15+@LCA?A(>aa:g3_f7=6=/;X6Tf&;,X:;/#P-.=NaVV-[PPWSR6
;DB8-25T8<BJ-PdGFY0=/<_bOJ,g^2K#Z17KO6E&PE2_S:^DX8@/Q:]K:.+Q.PX[
c+J1aM-C/ICZ+_#KaB>HV5<f(F;(T;beV,L:D8.2Ycc-J]CDO3]U=.E<(32QaaI>
BA2:[HMG(eD2RM>O2B&1)9O0-)[+OgNMHT<^IBBC9Q<KJ1L[=cR3:VBA6FB8LO+f
UHeg5+E\[>EO^XKZbG4f_KLSAf1Z,VK;a@f&bF0-D.Jfc2)LS6=A3BLf]-NXaM?;
T-?W4Vda8LX+9(e)BX^[UNC=UWdN[5>Va@YBB:aE+97]DWN-=bIg:0c4K/4L_G.A
gQP_S7:4U?&,-1:=>[00VH1F1eCJK3[a(B765<2S2B;>=D^RXOSd@H\T_8WDFM=_
.c)2c/@_#1De,^\KCCgJ5e1&D0>&T:?e^+Y6SA/)_@@e>7aIY@<Ue13I;Ya9c?3N
QTXAD^7gJa-I2-/f0&BKVM0&\SP:AHUFXF1=;&H,RbKJ1-fT0KX2=K1I:\LSaPV(
]WVG=P35H:/1_KM==OQC^J?+;;#@V:(B,b,7E^0/2L#>V@R30d[>5>V5&?CfKb7>
)e9<H;aSf/?23OLN+5KOPO5T:;XfF16FgBUW#Raf^N1\[1LgE:dB&[Q@Y@-\UfB0
GT961Z:G]gBWT=b._CgFZOVY(JQSaH4D?P2FD_P)fQIRE2ee>7fbZPR/3&@<R^PG
NUX=Dcf[3>B^SCV4N]THVRQ@fS#bITaBXF9E_:1gN_Ae:3^E62f)1NMH>.K4)Oe<
=3L2V3MaE0#c9/D4Haa&U_cN\I^Q+[09:.I72;DQM^@?(X>W@081W:S/J28G&WOA
/DPNbHZ@KOG1R___b&D8M(PS6@67HfE]U4ORd)&4E-Z]],(V,<fBTQVAL6&1L_O.
MU9B5\+J#4P/CV5ObC]&cd7JX@AC6T.903U8a^H9Z#cD9AIT[CD<H=ff,)0;HaP/
(SMg6:7E>gE6K)8c/b)Pf<d)1HQ&YgfVV3gf]S4c^](a&#-]#c_Ef;2]</89(;Y]
.dJ/\faI8Y#V?a6-fKES[VScGZ)EO9=O9QT@LYIGC+PP:96JJ\83>:/f/66Me4I2
.RL6UcCI--STP>J.PO2\Y@fQ?QfC-QCQ79>gQ-YfRQ-B<_Z<>#]I1A7L9dZ4PKE=
7<?-O,fFM]LZ_=3Z3R9Jg\FY-d:cOC?3RLcc,dR[d\d+FHP>^_J)HDU#0<MLDD]U
SUX3O^R@9:HLc7S4STO??Sb>&5G#R)6BE,G+a]13D:UZ^K.TC2],gf,7K)X77LGf
T3,ZL2.@Id).B/\0DM_P;dIR_7/D@5M#L5V]]84^b4&>MNU(@EH5BRb&J\ODZ+C.
^J7C>Pb@U-M#VKK-3@DZ>Z^8b-1MF6?&PQ/R#9[+,JUd8=O/Ye#.RLU1I]cZ/A?D
g_gUY&>?>]2IV6_C@MKG(L><b(Y=[AAW&U0gC4T;gO1OQ<G]7,.:E-bb97DN\6Pe
G52M>^9._]9fPM)TE1=P(473CE&O(cHQ(8]-&YaR.]RS5c=,gQ/Q@S_X-9a4)F[X
_J@3+RMS(>I<#A5E4=[_KT^5\^H3KfX]cb+VWHRN<AYIGB,_?WH6YfJH1f)4H<12
[#@(EcYH<@,0OV@R9R1F/G\+5.:#GVBf0a>VT_,g6]/.\EAV#VG1D\@OO+4cX.;_
5-3V^&W[0EC0=M\\J:RPEU19N2TcaHa_W;#_RXZ:9V3D^QZ^TSX&MaMGOJD\:M4H
2+FM6+H6[^,?G84^#G\bB0/X_SJ5;,K;5XXd)B=KU8PeIZ7I,QC^9GX8N3-UGS89
Mf_J6JFR&A>4dUAJZ&F->61&;8.b.>f34c)6D;H;5TC#\7.]+EVPH<3T<MP>JYRA
e95<bF9HeO8QP#__F_JaFaWP90b<3Qcd?F\P5U#,<YD,RC5PLG(VEBagf]+Z9^MB
O))@IA<&,T=YS].V/#_cE@0f4/>Z0bfQ1?N;20ff)\9TB6V.Eb;(DF-BD),];L>e
<Z/:H>PF)KQ,4Q?W+Vf(2g7AeEa:)JFbDZg8H<;S7)MW?3<AQO@52T,7;2g7C7&J
R<g]JRIX<V>JTN.aQ7eg&0HT[6GH8N.QW=2HN)OL2LH2B81#,\3eR?<g6\E&K>Q#
_^&R3TWVAM.VSSaSY&8fRbWTN2e:We:6O5-^(W-5,,._PNWD;VS^g1bH[)Ob2^1L
/LCW:0#5)]V_J5TEed+_8:1R<J&;/\ZA90GJV\4-afESCZ3KW\6[]bPV;a]4P[bb
C3FLTJQ&FQZQLegFF[ES6U_6+@K)YG^Xg\,2.4,eZ/aPZ=H.#^-ddJe)dDOY+d(6
5@L&c,NS+DgAWLNc@POL0V0;7MPU3H@1A,=Q-/eQ)[(^;gX:?:]P/9A6T=?P+=]J
F5##WTDFE2dTDD26]N7.@bBI;6D3:CCF1&6NGc_KXFg5O]#=;(;dATFUYb=I3ZNO
=QE+=SNE)?-a9/Z?1ENF@GI&RG>&+N[3\-L,S7bfgIB8DHUfH6IC95OH.+)T6(0+
;Y0DI[0LAUT6?\Id<W59e-HX8-@B;BF_[UZE>a98Y&X--/S8I/^G]-dU)UD((9\&
S#)[CDQ_g6+RMQ9]WBT:^QbL&_KY>6]gIIAFXO2PW:ZOM1,@C3YHJ0:\JDN@-RML
QP(c:fD-Zc)YE8#+#Gb)8g+[B]2ZaC>A<e0/OI#MbG^TNVQ2S7/M50aU2SVTgXO>
GPg4I+/.;6>&=T+C\X^WL4-TEHRQZ]f3A7#K3+/OfUd,Q^B[L>P/F4)P0/_)D4)#
L@9Ub@N6OIL#JgZP/_JX3)QX5@7MDYg/V80.HDg@f2[a493](PV5d])K4ZRKIe<)
=-)VZN4e:T595I;))VEVbM3@]FHUXV.K&B<.A<L(d+WTIR=;;O?7bd,c.V>E.0bA
(29]d14_#(QM.eO>:.Q<24CaQ6efd-^VEZY#Rf#&312:OAa&,KH:NA&5V0a_g;]1
RKMR30AZ-VV+@G=WFEM^[RM\N/.LN87;7K5+KKJH7=>(=[)#\]?91RB_^)Pe5U)N
Ub#.Rd=ZUa,@.)B0#.X\2?0MdOYFC+f[S=JU&]YWXL/EB+OA.IHXTAQ4P0^(=9+-
_XKTH,S6UKA4L1H5Ec?02gbQ#YH[DQDb(e@QeUWEM\V>]R]EI7N-C<LYg1)B:+(E
_,f]3Q<.:0]e0A/8McVcO;PM4D6VMNK2LU60B\ITR,<Y/3O^HedfSMFBO@E3EA>U
81;L7^99D]0TYUd;Q5XS#5=R.Q_NR7)R.R5S+V^^D20#]BBDObT_Q-7)ZY?D<2:0
Q/)E56Db.c;U;K9EG:#8fB2G,W\9e#Qg_#S:?K^^O\K2.X/X(a+@DO;\9\&@(776
,f_X,I2[Y,8JL<_Q<b3FB.DBL[Q<@Y?CZP\3\X&fC?#[+4&@Qc-:;M(O)^;Wc[B]
N@9@fA^HREV11:,3)dfS><H:b(QZ((+SgXe[g8Q:UfSW4IQ=:YPdJ]Q=H?O&#0Cd
&WF7-SC39fcfQW;97VOW?3^fNJ)MN59f<OCK:8C<3ICAFJ.P6B/</a=.D\._Da80
WZfKQH\IZO.E8;3cWWTH:\]_@KZcT,XB@21[WPCa2:0g(MKRMZL[TdW6/:d+]N_D
X=#K+INV.O4gT\78LGR9a.3R>PDIV?4b1VF4+)IWKK;OE13S^0Z@2-adVOTZ<He?
c3#-A4DE20<g,$
`endprotected
endmodule