/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2023 Autumn IC Design Laboratory 
Lab09: SystemVerilog Design and Verification 
File Name   : PATTERN.sv
Module Name : PATTERN
Release version : v1.0 (Release Date: Nov-2023)
Author : Jui-Huang Tsai (erictsai.10@nycu.edu.tw)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/

// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_BEV.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
g#LbA+b4\e+RL3SXKR5RLJ[7P\7S_)FB+<_M5#fJ[;UaMLOCEZNb,)2O6e[Z(P=N
LSX^BPU:-RB@9XGG[L(e#NE9fMbQ@<:CVQ[[84cU^M.R15)=M@]e#>@TP&(7N<E3
gE?EC./0R,aUGTP.2+L.Q]W[#[H,0fW19+@dY:AbdB8KaH_2Te?SZ:SV5R5#@N99
4L/J2RN^(GBM&X0D^0#0&XRbQ2cUcAa7;TR_WU1)fS5E[4(dfQ9XBOY4>N7Pb&T)
NWJZAB3_\.D3&]16F&,]OLW/<efgJC0K+>/&cCBFBX?M\C.[CH.31^3+Q;<EBB98
(5Y3gM_MEO;QWN;eVSS5).f8H\?RPY?=5#FEAbMHOD;J-g>.#8OG>1AFcc-9T<-\
LV3L3fgCJZ3MC]I.AYH,I,SBIK?N#4E7P;c>>1]659b6_@d.daT1#])RLIJd^KKa
(6YB-^f4XJ4J928b)N&N?RYU[+#M.aDMD<<I;;&Q7&P],dA/F;d3^,.5V&GTSEH4
>X3Tc]97I(BKF.02Q?AfN1N83\P<A;HaVA>e.DKOGQD>a3U1ZYbMeTKggV4U_?)e
A9;23#+aFdgY6QfFL\);L&f#M7F-ND40DZIHKTgF&<TOe#COEfO\SedAc(:[7NAD
&b)VJgF8:8-Z+]+K#A(D9a8;LZ7#A\YRcP[V+9N/AfaC2Q:g4VW8&E?[,5495@F<
NCb24-c:[3RXJ<b@E^TY#@+JCOU7PbeOY1bIUP-ARK4fCG0_e+&E@WgZ,VZK-aWQ
-(W^R&-1R.@I][WJdPBOdR=<B-R)1W1F7U72:K<(_(:_7f:U:\VL5:;DR:eI_XHZ
#T#4<56Af.[7X/@02-]-X^dCM+0;)5]HfLD8/d8BAeb1,f=NH_^aV8N50FK>4<dM
L]MXG5M7OZ0Tg8]P7/fb5LT0bD)XfRcFR,I@S5>[=1:bb].JJN<<b<AZ5LQJ)WSI
JSA_=)H9SC?A:N+=/RP+LXeLgN&8cJN>\0#9^6TF0:,f/577\4]L&LdP8I,XC_>V
M@MEeSIJ[U&E&O.&0@G9GcdYc.-eH#VePEX1,4XB/VbPFA?(?9L/D(S^1AB(?9GU
K#02((I(f<UgVP^<&AabDC,N]VTET5Q80.VdR/UJ_JA:F5PDWWVd,6cXVU>W?XRa
H,b?53E4#J2I@2DM,TT(41.2/CB-\B2X<-b21;U;G4&<:X\&N\I=c_C=]VPJ@3LS
X2-\7GWX@_3XRV).3H;<9WNBO1,MM_gX9AcFZ\4X,bg98T7Ie1N\e3d3=/B0CPQJ
W76#.B@\6aaFff4(H[,&fM_>&B;GTWW2e0N;,@aZ>0M=(57JJ#Gb_N:5SU#.MV+H
9)1T@9aZTF\[^^Q;H@M7EC>FKf>[H4aZKNYS3/A@WPN#&g8.0VFdG9(JIF(_Y8-)
A5]S.eS,/(L,fF?DE?FM2fYZ:]gLG?7)a&aL8\A25+LV9f<G+F^#N@+69ST/QVBX
3.?g[g[R:3O-Mb_J98YH<OX,\I_O8P<V,@NFJX#.0WF+e^^cEX5/J0(HH6XL_1c#
T?f-:;&@E+U)C)?Y58A.,Y-fgAWIMV?1IGYB@_B+@86S(;\>Q7SPT&D6:<;3\PU2
/GHfQM7?a^c21eDU;1:C4+:9ZbF96O&=VL//8O;D5SEDAFWQSga2N2dZ,RGS@5DH
eFJacLGFW0VRRMBMGb8;ID\c]MH?(3N]5J8:A.FUV<3^XgQ]X<NEX<J)@Y4fY\X@
DYW&d(c:6?7d4RH\L(,a#5U2QZcM:#6B+,?=&:?<S/.IUVLNXE03VWEc6-V_\UZ0
1adAg-WfDZV]Y?3aY0bdBUL13[U\@=4/L;9dWHNKA0,\DN4(+(TeEK\&5Fa3MOD=
6ZF^R-2g+YD(eES==A-KAC3>f5]/BU]XcK6cOLMQ&]/55b_?D-8SfBLQ:RX&g(A_
BRKR9AN^_[UR@<=XA<?Y8I>de+2Z.0Qb<W>K)eF2,^_H2F#MD9&FNON)&2R#QVN2
ea[1X@)P\R55PS;)N5M99WNN/JW=M58N-W_)^3DQMES9GQ@a1>/XVDYaKd+95JV.
&S,edd0gfaNW,Tab/V=X?1fWPJ2=SfM4M&9+UAg?1d#4P-gOd8gg977&[>P]&O[^
>A9FJ(cOG4LID+HLMQ[?IUF/GBPFI2MZW,=U-X;DEbOO17=b9^3M/bDW[QZ;c#C8
HZ0#C_UEHSD0+SJES.<DgRAG9:1dV&-N:N&[0SN+e@U;=,_<1;-8(H1>R(9)_.NX
eNc_E4+(OE+,\fN<V9P?G2N=7b+?a\1(<D(G5Z2\/S;M9E<.Y):(T@A6WdO8)[A[
SHR48[<=1.AE?UQTTW\GEELIHTg/&L/,deZ1[?_1fB()IK4dKTKK8RWVA]E>_?N/
bN_bAOC(@O2aC+R5f(QY@?3R),@#/-:OaE/,R/e3V3&L-@SAANV=F,T],bUP9c^&
4CVFH6P:-<>3IBAgcd2HcGI3PX&FI?L,88ge)Fc43Y0JXYUG^RCS=<4NMRAfL,9M
H6(X:WaQLYL[f;SH>eWE6F8_@bX1ZA:5NI/dLP9C(I0J(MD(<)I5XK^E\O1CFH@K
Q[&cM2=S=Q4(RGNU=(=,L8Bd=;--[-/H#M5;.T)bB39:Zc?E]66\B8DgEA5,P]RR
._MP4D/Ab]&A1BP8f8.8+R(D<[B<\TUW.5Re0Z#X#gKV,Q@;50^e=\@O#?BRGZOA
J_cAMO>W1eQ@+_>dBN>eZ0&12276,&)Y97YBY&>d455Q&=CcN\D.BeOGTK;Q()BH
YH\_BNHQ1,BMW,gMR[D:4&NIP@5>;LR(Va.;3.fA+0Ae2.64=R^S4.6GWT_B(V0W
679:,&1PJF(3,B,_3LNO]S5^bC.,;A0g3H-,+@D7T#AcD71R)GfH3Q4-&CC-c\&0
B+.?=<6BEG;^KI?;\R>KRNgC90\4fY3Z03#?bEJ0]a]^a/++(U,=M:-&)HZ:A+9g
->G1B81Z[d2^[4W-#]TYe6e(;^MSd;[<eCCV&<)D@g\WARZH>e;GP,Ad5&YJ:;SH
/#OD8)Z#)/^)MST7c[YJMS>7+F)G8X(8)NfB9,\C>R-[2>L_VL<?;)Q>U<TVd1^]
e-KFGCW,-P8^2e4+Xceaf6ZgZd+5OU^L&O6_0E\8B)D9?M_Vcd,4;>e)/P=B\D<C
WS2c_CC)\_)Cg?eE#0NDFSdZS(3C3,:gS(&aM?XYK;b5d>P^RXVV(@b<A5YIGY@a
Y]fE+Z&BI5gbC9LE#4VD(#EP#R[G).(D9EW[L98Z,UD=Mb7P.E2SVNC>>-RYeW6Z
#G:BD.;D?-@R[Ad^2bKHc\dMObAV-0;INB/,U3X.L828[7SM0]6W]A/;c,^2NT&/
?-&UU+cT=;[5TFacV+2LT0V,Le7QO8@)YG(>ddREKKE3>8W^H1NVSCgaKaC-WH=b
-IFBc,)D[V):dgZ-I:+ODa5/SJ&1HYKQD?_N?=&[T7_d7ICLVaM&)U^2TQ(Y+6<(
5DGeCOUIZ4O_LG\B956<G@5(,V-YOA+GR;0GSY8TX1K><Ea.-Q0\=,Z@5/[CB5A-
S5Y3\[<2g9+@9.;(4^7)Y5f]/5e2#Z)3-F:EO?T/@GTPGb.KL2YeKGBeV\Dg81<X
gaKVO?6R9BJ;f,9bg[b;d6/+8f9d1=QGf]e-A=N7gZ0LPZ4O_cPf5&P^(aSbb19O
D?O7_14c\&)Pg2V),gQVc>>>8]Vg6ff8U(4D.ADT?a.[dfM0YDDeI[NENZ+KD&R#
STACEP8>@X.)2S.Ng+8(__[K=&)E=&M211G]_XYEG=VJK3[TKW_X,:P/XK;1cY:Y
VL4#T)V@Jb55GfI_U(B6+JU_B;,&.Qa^,bPY>@=INZG@299();=H(]Lg7A[OCf0=
a\F#8K[b&3V+7:aeM<[Xb([Q70UULVa0G&17<_>X09XN7)PJ)/.2KCN>?G4/.&&[
SZZCM?Z@7c-#]2,.9W]eW7d4eD1U@>B7:PS&bU+fa#[2H^cUB>94AKH:5OB\K/U\
E3TLc5eT&8KaagOLIZH]+A^649_NW;2XP2g,(UaSY1Y<]JO\]0+TOKg^/GG7MS&/
-P>=C_S]_@2)<Sf[NWH4(#KcMdE&L5a]7VI)[8U@ZRIEX@.>47_B/WQMQ/2Vce@^
WP-Z4#Q(fceB0e#bUNC_CZ0)TXGG03a3,=?ZIU2FZeVLJ1bFX/B]K;/EM>d.Wd,-
C5Q=IF_@>T?L0VD:V&Q[CG]MXO,=6Z5[?)-CgeTMO.c/5T-?K9OBN691#-43;@=+
3\>>86/D^Z=6]43,eJTg0,56Eb3C?#2#ZZ)=]XgeO/3a^C:00CfNQ-.3Z2DPaN@X
9[H^/MG=6APH\PS-@>VHM-1YbC_Pb,]6VOE&UbPHYdaV?86-@-=H@8RAFLX?_V+P
#g5+Ve>E[E&>S\Z;DIU^@eKL_7GR#b5RNF4LX6)H/]FJ47bcK[_\:FL:0_DHY4S4
<(9gG#<C/2c+1X1V.PD>.c9O,gD@&ecHJ-UfI:&9)(ZSU9ReSg)O6YB2eL,/)G]-
f#=@T)a;0QW8Tc+Q)AY-^P1SML)5f<fUVVf]EHV+3LQ.A@@/8QN>2+TN1.0c</(V
[Q&U0,N6aaAXDGH7Tf/_HdWERGA:Fc51+A^6I+fAcV]-U:C3=>b?V3=^8eVOZg\E
IgJYd)P&0/P8M[>.f/\T4g@FV6cQ2#:_#(_WaHL-12V\Y/>#E_FO,9f,IR+b)U@<
(WQQLL6Tc.NLf=?&F46[,A\B#;RQ:^#10]DbH:)Id1HW+;)(,-FXTd2L@MCB2LM1
<XO(,A+,<e+?U1#BB?-fY>@Q]-e?Y/8.9g0R;82(2I>2/+BWa_J,?#]FF5#1F]9#
:LT#1=<YI88g]O]-<gd:fD6VHM=GHAQVO,S(gb8CfNN?C3WS2#W1=a^U@d/dOG0:
SUgTI,Md>-0P3Pg.8H,LY;R4g=L.>fO#dK_#<0AJOUS?,f#E3[<OAcB,-]CbDQ2+
cHN&81e175IB_78UgW7A.VId@9@C65@\Mf>>GP&M3^:+;.+;X_d[-;[:N^<_aQ[f
4<39.P6#.QVG4gK,=#MEJ-.g0M)PIST?U#3^8R?H99>=LCQggc)f09=CVe,[)@O+
9M^DI,4^+WHQaR^d_;0TdV\O>5M9cPFL6gZM&L;3R9X?gA3]A+PY40FO-A/ca8Se
/&C)_LR;X91@2)NLRf;LMg,X[K;+Edb^/OBd_)I<9/-F//2XOEW-gQZ[#DTGOP,7
=LW;WLJI-&]+^c1R<fRG,#TZd[deXC^M?3CEWFG8H2-1a27U2]cfHIaVO&@Sgb?_
XSU@<D+CS&IWYc]JbIB6_5QfTRP?1J_:+0+AOKbN@R-/YB^BDdaVUb8L3W(AK+\B
ZS^6T3_EO:OB6(99O4\@]2JI(fb;JL1ccZc\e6eFARgZOD[&Y?ACf=J&AV1]#QEK
H,.&S0gL=?f[D#WI>J[,.:O+S#GZ-UL&eP47]0N73/^NHLXXc29P3bO#W28VX7,9
C)V./fVFL5T+=OfA5J?O@7GcD<<@abKOXS#gfW\YD(X5>/XgEdF4)5,1GgH#^M5f
S_fJ>&?EK7(dGG6GE3b-TPQ@^]L^C<[D6=/DB57[P,#(ag9ePP5#S,eHe+@3^:\.
Z#ME3S8#1K<X@OFE728J7+O#J?\^cf4&.QQ+E\f-L?2R#(V3.f<S2I1bE]M+1DPR
8bHFB2B\6F-.V5((0B#1(<4W:^QOR<2B@IUNRKeB/.FYc@;\#,+53;&6<Y/Y/7Ye
PI(5:&MH>dDG88@DIXbJXfU.ZKccbUD&DcMbcQ^5\;U[)/LAZ\_3^fLZ+cWgJCHA
QKMWe&QXLO77M4B.GC0CKDM6^6de#S-dA6(8>NV:\8A6(GP-]c,;^7+VIV6SW>/M
:IBIKV:B,64bW_;7Le:^KH=U7Q:70Wc_.RC/-T4\5Da7)MGRU(Ma]<97G1O?JA1K
Ed1K^=JPa9DS=8QW4Re-]5]_L.30(JOI:edB?DRS^WT_T+6E+LG4<0UG-FGH,&N+
G[cD3\@L_aHf29_Y:]bBEL9bS<X2aL@X,4R+B2QO_@ISc5V]?LR9bF95aX3EA&ZQ
0dJX]PFK[(>?0H#WcK&BNe-M<U\Yg.6K,F-(d3E:O=+e+7gY^=@)NfZFUeZFb3<5
3U/)UW]bb_6egOHfbc=0+/:2[K19Lf@,PDe^JBb\2)EV7/deVQJ=STMd35(BF\@^
cH5CA7/<-U:>2bD157[DNe<e0c@4=1=eO+Ia</55-A?.Bge9OGe[eWBXF#VH7)eV
bKXUDW+9[?7S3WEaBd</f:05UIb=fgM(Hc[V,6(X,@6NEUM4TCL9]:@/bB]1G<;R
;PHC\5;]@GF07HSXADKDYWU^^?e)>)[(<I#g#((Rga,I;J<#aV:?Ic[C918g0.8[
(b^5ebBW#6:=WLH8;5XDIPJFcH:4d<=MK<:H7>-dc89&T)ZAFU\GF.,bM0L+-0g8
+MT-#@U/LQDFH&#5FbW]a2-.4F>]_bZAG?8dWHJRV6g(\gbKF57(.>2:PZX((c84
+QDA4VfOOT\1:ZNLT8=XA]I-QY@YI7a9e[gBYG)9.#_K?X7I_3A<P.4LADRbgK\X
<=?.^#a6I?0V/,#QJ43WRW&(#b0BM-WM.8H)F,VNCZOMZ)HWP]I-DG&bHf=eB7=4
f&RHK;V.;>ZCE>&K&e?d+=C&G)G,E\U,NB4\&4ag#N#.\N?<9(BP,bWEUNfFbOaY
c;44)F.e#F#gKbb3B#7,_^JBA;_HNAeD](J2f^a#,WG<S]UEdf>2_ZY+LG_.>&@H
@fR#AFA>+[c(e#.ER+KIAF9T=/.A=?0=F=TR,JD110D[@VP.LVb2I,FgB16Q1NPL
K78Q30aUFVA]-FR,b9@b(6Zb[JYZFA9.3E1aE8cLM),Y1TV,^IK?18g_FFM9=SCK
Yg3]8P?#I?JY6?W/S09WC<9:N#IDEVa@#(_7BC9g]dd_f0&6/FMHHMM<ZL];4b,V
beW[fWUM/e),>;@2PZPB+90fK1-aaV1<X@6O@/:TS<SQ,>g#0U+CI\<EUU,b?:+Z
Z;7f\M&G5cbT+3,9&(d;-.DM0137:.:LT@2V\NM\>dL,]WCeNC[60AEe12e[;cV,
R9#[b:6=C;DF2L4JCGgL[SQ&49D-7b,[JL.1K8.57/H3]]P2<;+-TPGB1H_OKBG6
IC.FY6]7SZ:aI>XI/@^X&+VP^g;/]+?)1(J[Kb<DM<]+c,eYf/[ZP2@>bME-NXUF
_Eb/+X>GOBb@@PJ3<W>RBFMB_PT+aY?Mc;7)(]?aZ#U0[bA6Y9Pf5BQS:U&68:L?
C^PO8d1[cG7-D\60Q\96=09T:G==0RP(Z9(5P_gT5531;K#EWF&e9a8O[J&]#Z^>
Jf4gY8;IE.C_T;f\<eR^X;\SZS@8]62b^F<cN1gBB^Qc.\>,E4RP594_cA-2E.,d
9+13>(NgK1Y@QXU8Ha)V-+U,e76(SVd@-R&gN19E5F&Me_;:(1Q?NaVUJ<4+,&V9
6ScaK=U7.U>:F@.YD_^_7Z2:W^;g3)74?,X9d/>Sb5LaEB2WCTUK[\-6&fL<cKYD
J-0.>^(cU6_+RJJ\O.9OVR[R:X]0f,=D8)e3QB#S)7J:X0XZ,Ta/2e(Y?IX=X+F@
AF_+8Wd>GJYS9)b4(F[)W&GbaTK6Q1@a?^^L#aXNFZ10W80[AKNB-X^b(6\>fB6I
FcX@:ZAD7T)d2Icfg#J:\6V(LE(W\eN/&2e34,@=W/b7+(a\4g/FXI7Xe>9J&&>F
)9RKS)ENBLZKTO#[#)U,V;:R[()M&RV9H3Cf<8KYGcUNZ+).U@#R+f;1Z0fWaSEg
>^5]WK:7_b8[@_4F9g[V#b#8__UMg?1ZV75.]6X?M9aAW(La2DHc+eMBbI1B]M0P
f.ef[a=VK4DEIVIS3<G.WSZ>G\cc\AH1f#4^DK5&2V0:VO49f?6HgHdPYbEDIEM0
c8d1-OJ2JC7Sb=Q8YN<Ge538]]+/_P?L6dBW5_U]>9T?(M#:7fXXX#&K^;fe939I
C)A];]ZT+S0+MLRFAXCBF6\g#Ed]PN>J[_-L0;^0AX+fFc>LcQ>-ITHD3NK6)HNg
N]#C7][-)TQGD<=;DZd[J(GPXb[L^G?X/eW:1.La_R];B)4(4OBe>(E;8V0K-P<.
dM;F9=b4>eT-f/8Z+C&[B8bB]L(@LX^Y_EV(dSOcTIXM=5e<?[3)?;6VG#_P(/NR
dWGU)LVd6HWP#,)<&\G2W;OT@b)6-<V^@][NAI)8;b\CE1FP>LSITTJ=K_,ZWf@B
W-)WT2_75deF-/ORNR-YZ>GY0c6Y8N0F)X5<M<W>]9=#PS;^TD5g_3YDad,N&S&S
]/gfV,=&YQI,[H;>+=I8_05,-K68RSV<;gf7a7a-_2@^-<3]<F9ZQ#Bd.UOa>KbJ
7e-)_c&G=XfYA:(^3POR-ee0(/@/&YTHFeJR_&JD=(;]9ZHM,KD5fLa^,#VRPJRC
.IIGSK[eHW+K):bEBL=SbSW6Q6:^NC9Rd#^/J]38S7eSOATF.F+;b0?LfV4FNDSW
<dag,ggFTHa#6(MF>Y7^[f6:AXQ]>Y=fIS0YVD,1gB2b1X^O<R?gFcOK0Z\c+&2U
>.HLGJ23\1UbO;f2A/3P/K)TYd1O<?]/8gb:eAXK]6cFJdOCE^12US@,USg+5V0C
KLc.RET,;;4]N1?G:#-7.Bd>4.S]7^JQJ\8?5K@-_-N>V&OH=JE<6L[Gf9LXUXJB
/JNVB,4NS>3aG/FT#)FIA#g^Off]eQ;P\gePIET_@[#d-@.\HX-^,G^[7XTSEMQ@
eN1SOK#dLL6#4bN1#5:cHX?JR<F(T&D:#_>R)Eb<HK[Le)A;[097,6(VXKH#YBQH
J1fT;DGJJ-HY;@Y[Y]fAII4d91(Q@ff/278T]9).ZZ_2O4QA<ZX<6OeX0dfOcX+H
Nd6(52Y;LTcBLYe;I.B0.b8SBe@IX^,^@eXd)0L>@<H_Q?LZXBb-5F2=KI]f4DV/
,54Z[E)ENR>f/d6^=C85VR66(E3I_ZK\:SQ>4?^8/1Wa5R<#P2A,P1?dg5N71MdP
+.bKR,9Cb+LT&&U579QO&#R>Q;gOA=O3:_LZXQYNe5V:8]8\S(C7/7TKRZD\V);0
/+IIK]59O(RDP1SBa@TP]F_ZXPUTR;@9(O8W2#F#M@P56[GQ0:KRPW[;5=D8UJ^Y
eb@F+,SKX\6eZ1Q+I_=J:NEP8OANUM3VYQeg.9Z#37(8O\R&<X;ae+S7+dM(bLH<
(UNf@(g>)gPUET[=,\7;D18USK_B]DW34.YG;8?Tf6JX(/CG&E/T;3HL6P_<3.N(
1)+&:E1ag0E7e?^LC>+Xe(41D3DS;OC+gCU?=MC.RDFC7e-\#<^5(7ad187/a\7&
3?0YS]G=H?-AM,9,P8NIc,-+4_VaJ).fAS3MgDD1&UZFWeAS]b)H;bca;I(\Ze;N
HEW(SDCRLEgZN0U\P.Xdb2>J\S,UU(f.H>3#g(]:B5C6>>ZR#74&)+2Z(eXKILf<
=_8CND8@F=)Z\0INWCcR=K[[YGY,:d7G5CPB/8Mb&)4P6DN@6-P@,(),#((DHJN<
J7^T_^5P>MF?7bJ-cNaOEYHG1]gSNT]<Y/)&1IBFeb7M2Z7]F,[L.[[0[@AU--V0
=8D]HZ6B@V4cfPSRPfeACWSb:_>GG/f+(&]P[4L].<14.TYMBM<>B:20f>K;O/K@
SVIe#;W>Y<:P4F425OG6NTT-_YEf2O,7M_g9X\R\P47:VGGIc5AWf--33\2SQ&4#
YSaOUecX4<&GaON#/K.B38H+b^2A>fF4PCQ0YfVPKTe9=<0b:>HB4/U4HW8,a(PI
B:K.[L#D8NdN[F.dTU6fKYJ9Y_Q\^cPU)TKR(OX^QJ<)H]>D2Q48A3dbTQY7<R-E
4?YO_>+[ZQa.NRB@25Qdg4I2MQ_1Ef=@F-D)U^3S)@#;M2\4Ye:cJeJH9HE?e3)6
a+^@0+CeT8U.==;eaCFCBXfG3U_7X)L<+EE8[M1g-J,>P+^@(P0O&O&3@fY>PHRV
RV#>Z/V8b)OH1SKa-@,0TOBC4Gc[>,P4Wa//<F)d;Vf4^e96&cIKZ(;c2>Z;>=EY
D?ggG#^gI(AA&)KQR9&-6?7?XC18U\K6cc9W^2g[(3KbXIf(=JgUT+_?[)HV&Q=G
CJ1ZGCJ_69G=C7fa1POcFAC@IK@WV1J4aIHH)_A>7.0\;/E#]G634cYLL>>b/e4d
E.K()Pa5?\00,OaRISY8^<DD6Z,<X]4/1T4ea)9C9&WWU;9[0Z(gKa4,K0\0?-X6
3VPI7TYD844Q+/8_>Jd+L_/dbe6^YDU;)NI.3>]7#V5d0#02NOa@@eXgD;6->0KQ
99+,JFEB(\?8Y\E=62-d@<[F&Uc[+gTM74<f^4__WcGFF<0F0P1Ng]G[&()KSI?9
+/1&22bMX@;CLJ;W#IZ\7@^f=+YO[b&#\?Lg24-e8eVa[Eb[^d)g:F=I9(LV2Z7>
I^S:RSQ4LS&>RAWD1,]&XC?TfO-QSfOOQ+/MF[Pb[X.4V]TK]KU1<6Ue\e/K;AK+
UWX593@CVe4@5S:.dLb=OfU[);Z.bMQK;R_4+8>F8V>MWbcafG7+e+aA]19;NfKF
?JA=&?SMa299EW^7ae=\<)?g4E=DX,POe@1>Pf?;G2e#^-4>(<8?ODI4>M(V;;:;
MQdO,L7aKPf5\#1/5?8^]794PNXcQKd6ccJB-_77Ibb6B39&eB^Hc=K=c3^7^>cF
92Gd?D:TafbLdGN2C(3\QBCTPe[,^8SGGI/Ae6cA[\XZIKWE3^W4baG]@;=f&9eg
1<5GW4Jc6KfUQOS-U;JM1B4(b[G)gXJf)Qcd1f(7YTcGF=23XC3_gIdB>>_#<I@S
J+(ff=V2O-#-GRf1;c?K9K+=-R=<N;AdV9+SS5LI1?T?6T?cM#-M@J<9?U[;Y&0B
&NY6\5.eA1#)e>SV,AN8N0e00Xb7@->?cVAB1-5fC0.bbgKL6)cV;+MK<A(.^]GU
@Z1BaZRd59FM9K7]XVDJXb.U_c2SYfO@fL4ABI7BQ[5=#eWIODK.V#GD@YN0/OY,
-/]aU:P8@7b.OZ>\9W(a@83e/0I\FJ0_#3_<+@&5eU5YHI0da;::GZeP)EE=2=E1
GJXc+6EG5H(8?AWS)J:RJ(SP2Xb,(_?877eO7c?EN+g+D:R]/gP1P0&4E6RR2#,M
aQSCJPQT8:&Y=3TD;=-P6N.=[J,6]4G#H^Y7@g\0CFN0ZWaQ3Ud&TD45/Z,&P6ZZ
O6+,=<WNeK4cJ(eH]^S@;8L<<UBX-U=Qc(BO#[K^M18/@MfF\@\QR[>dD#_N:4/2
A8D#OZP]@-7B80WU+M65[-BA((/3gM/8I253GJ(.]fL&8Y#P7^)_dU0Gf2/0L;YZ
O7#GC[f5cDd_O+(+SMX^,\D,/5)871UUc(-7-1ZY.R6&XQEYRObU^0^K>^</M1P[
gRPf)8QMVT@4cg1SVacHfFc;?+_U0V._T:XSI5DICLGS<C;))ICIJ^cD7=aW=ZSZ
R)_=XK0\2\Eb[0IKKSA2QfVD2,#9;?BZ-HZNEG5:DPBM1U=@#aC2.g5RIMW[TC+&
ML<OJ#WJY.(Vb]ecGba0W;&89U=IIR[902\2=>3U4[VB)EF51bZN2Eb@PYIe,A)8
,2IbYUJ:SI(\[U6KgK3M+_[Q1YJXa[E?>WMM3@H..MYR&GVf05L]Eb(EgMF&JQSX
]G?FD_g@JDQA+;A/B,6^LNeYF6OAJa[3V(,V68MC-Y=@eVgK.EYgRX4[1ZHOB9_3
eWEGI>0@QBE5U3]7[[J[97?71-I4Y,A7)-:426[?K^M?JJ/+M.Ya0&??@EZfU()P
^LL4G@gc1#B#<:G]M&3(#&IA:>4440-3)7>b;B=;/V7;L?SY5YO=Q8D.XeIK(2:=
#N<?Z6Aa]4H/d].X,&eC<bec0NNVRfB/TQ4S0?eKHC\82TaeYYaS3N/P?H=CgAc,
K)^WWMEXO5TKCL:]N[N],bHEEeH_GTEEFT=#8;;F??@2eRLcEWQV3V3H5Q1bH-VF
Lg1E@K]).F#9S==5H0G]cbaPTH,DdMN_4I]PSD=VI5d9IcNS^7B5=GK7\YU^A6>5
<-F+)^4)O&69Z+70MdJgC@R.-7A4@UfX;A&U3\A:G4<-D?>&dfb=/04I@^P[g2V)
N,FB))g<+TbJPNA4BgV[J((?UTF>2UdddZ3,&PK]2XF+J,N(7gPC7Z^^86aJ>d&R
98-NEDF>;2DH?3H[(-NE[MIHNP]NSLF7O)]0()>#]&f-ZX<G]01-ZG0O+)8O#5gH
_c_LIdCgA?dbAPF(FPg/9IE0X>e-6/@GX4Y.HGOG_.DgJ>&3:;A=YAU;,c/Z.Q3[
]8[UTJEAQS>@b0Ye6NeV^XMgYcZF1(OF#);N\Qa_e^84gM1<F<FWP.7XXGKF[&I1
Ra7Q#gW2Mg3[URd;@NQaPIRB2e@J=Y0_F@KPEY@;I9DfVR7KRVP-&QR_54Z7U7^\
7L9QX/(6C_&L85V&)8WE+)ZC^?MRY.UZ[0L1Y_L4GZA4Qf2L:QQg5310CM^W]P1?
QIEg6@CP<O7,C62e/4g<fIT,a&#<-LW2FeF5O1a+B<S5>\EY[>[P9THAVXU^7BLa
:2)-a&ZGL.DEG3.I+S0<J/)ASL.:4@1N2K7JY?WMN0A0G1\>&F+O]LIXCN&CIf/?
7Ad5A92H#@^O_+bBV,VgE)/S=eLg\gSf+IW#Pc<Cgc8A>Z/]eNV]@3YgAKLSDUJ6
fY>fdN<d=1\U]8f0633ac^ACQ@)Z>TNa<\^cS>2&[:-)R4bRQ,XaV,&Y[K)-35L>
(gcbYP>L/ZHdMXg7L/^141I8+LGcVZ2Z,BLV8W3MF4Z.?:4-X(]VPMPLDS3ab+@)
=V9&/#\(-7E\<c,58GKH5fW2EEFN3<E=6M[KH>BP#FLOW@<2O@DdH[fg[DB+JKTd
G?2F05KG7I[S^)?2#)A.XgK>WbgHI_g:eX(MZPM6[fc]^-IE3)3Y.ZK9<9M/9,=.
QZgegKFH::4K>JU5/b_AT3(>N56dJO6[_@BfV:VVJDVDEIO6P?5XK-fab9FLUZOd
F[H>4YLC:2AL9:;)2^8AIH8e2[1)T7LVgXAK:0cZ-EO5g;9.&I771S[eA4Ae_B-g
JgGA20Z>Y\cN5_.E\aLbZ/6MeFD@(79U-9@aP]8-JQ[cQVc1Z/J>1S?b)+d^;KK2
M<-gd[)a,c\-=OG;8/<-E<eXDWXWbFd6)5GOG887@/WB.,-JY(+#2fP>L,C6?.NT
CA<G6FDM<;e8[+GT=5AaC)a7GSW1\SXHJ;-X(>EH]VH;]7XFETM:1:>E9cFYW+DM
3M@3S1XbTB_-^G=1L\_T2V2a:+G6^6+0B5U\O/1DE=BV3FaJLgcSFKO[MK:RKC]?
>N?Ff5+NY>F+d)d=,FAS4e#(N12EZWfbd[/:\2U?)]JfKL@];BO>R^SVT-Ma>F:0
IbQSP95;0VLb=@KUa^(WQ/&YgNK=.?).FA:9Z7c^A_QQKX1EHO3LaJ7+#51HM6a<
FTT];7=E66@d5?/6#65N(BY\PFHE\>WQ0Rb&HQW@YBRP>+DDN]c;Q&QK?Xc^QN)_
cdBf0XF&Vc;NefCWDC4^&V1?3C-TGRN3Zf[Lg4ff=07)J[TI8.+>(9@XW,[YT4DM
F(BOR()g_JSEUT_aZeSLS0?=<@H8Q1UgV?aZL@CYZC^Ma-,f>NM=f:a((6&bMN^B
9U2=R,<&6N,[GMM:#IZKdgW.\H>G?QB5X.\_AWJY;E5AVPTXfL411)VFCbDK7&cU
G:gebZ&;(@SHXINE@]^=W\?aT[/?(,eUWF=;.^(ULN40KcBd/NDKIf.XL9b(#S-#
_3b_WW&\VX(;bg],b^&#f[e?X?#f6]5&7Y:2UbKM=<#ZbPG6D=255dSXg(T:XH^O
P63.@7XQLMWH4]HW2G?&_N.SfEL6I8?,RNI#]C>BR?6<_35SHe893S?P+G-485\:
_PG#R;/:>;AgEU\1[YWKf3PD?=6GFbg,<Zb[X33_0J80&>;5U]5/7^?Z=Bcc]IFg
54/:CD=\>MX@.f)PG\D_<BWQZO5/CDgOC/.N9;?.Z&7A+-B;\d<[:&dAJ5F2/2T@
5aL<0[Y)g:e_U\/8#,(DNWBR_fNIV)G+(G;^-1F;e(6>GZRBG,IfaIU\,eDWRAX;
)XFQ(LBdEg+aW[cb465bNDB;K[:.S(gDg/BC0)_08&/N9;6?OLR5^:S+JEW@6Y6b
FGK^fE\1VFD(S,3=C.V,-(V3PP]6ZcLg@U6&DMZB<1PMUAHZ/d94\>dXB/Z<#-Ug
ZW^56g88>Mg-J8aNb.F0O?9&0YB-\JPA+beJK@\S,8@?4-USXVJ/;Q@gB^R_.&<Z
6KL/\/UI?73/Y[G&-R/=80BMV#J2#MAEL?W&#JNU#F>&:YI3X&5U=C@E8JP\N>F4
<[_0G@_@3B&H1c1NF(,9>=RPK:,8A<K7G,Y>6I\UdH=H?#E9Z9-Y@W>6&Xg+GA48
627P;e>(cB[V@(=XagC020:QNc]e3CU&+3;^I</[Ub><96-e#9\(Z1S<BLWe@KC4
R_4@<)RIH]ZB&_\;&QaD4d+=1Kg_eN.d7DWdLU2[._2_F5;QW:W)USL)/dAeAA#U
BU)A>@c]P@U^_30(QW7+\0&&O>G7ILTgX>(Q?ffbcR(1K0#28OFH2H8Ab+[LO4:1
@W8?K[T>SB,SK:2WS)RdM(FFgW/AEJ#:FI/T)RCM_APeU=:^T@UUPMG[2PWN4[Uc
-B#XgNJK;MGA^W-R28RZT-X^#MFRL@,d\)?P+9^[#7aF.3U1L/\>2I&<,.#26+?,
DBI1)T<@@=64e(2&5^E<.PEL;OH&S2[&Sb0bZMA(CUgbN?>GDB;Vg-U<U27W:AIR
L8C(^OXeIfU;f>6;.-];:O(/][g:ZQFec?=A.N,Tf;S.>^@^:D=@H])=P?K/eP^/
9[+O<7-b,aYTN4P];(0b:9B8M>UEB1Z2T;e]^\+#.J\?<7-90MF-AHG,6>)ZI),.
OA,S#0/2Hg8+KX.NY:Kc5#&;:0+/Fa0a5Wb7b;?[5?@6-C;N)78gUe]IE6Z7+F4K
.S7#-6R&S)e,L,Z[+JZMG34bW0BJCKBSFA#N,::C._[W,MgST=[R77_6.URS,#.A
P-]B=UD>#CR\?&(GeJge+))]cK;Y&S)VD<T^\E&0@H7;gA4JgN^5\g=LL2]YGW?B
.9-(L+@^;=]L6Z_5EMA/9DH<f2D/K+#_:C)AB8-+=BS8T_f(Cc5.a#0F+Y4)R<SW
g;FUU(#EWbAf,FbGP\U<]<W1M5aQf\88^/?IV6_5a&#,c^4E,\8)9)Hc8cVb)8].
)2(<=Z>AS3WYH#N90V^+4)c:M4;W/Q:.=NLN]R8a==.g)JLI#)Zf=3S)@4aEg;U.
a5@W?(=[If@V2-;+627g<9SL_MAcVP4L459XRYS6@_MLgJG(_K+af<=<LeXFR)T&
=fQS&6,D<&U_gL=f0U-d&9C_>XGJYP[b5:>A@9]-B0Q\(]O0g3T)44[ZYT,0ELP6
V?SIJAB/.6PM>7^2f[d4aEgX;.IOIZ0YT,Rb,[gYD=SUAC711(>X(#gUaCI&/Gg=
,:UMI^Z/d?CV;YHX4O1eRA+;P\8X&6(D+JC02b8]Y(W\CDCFM&,;JBc@fbb,>-\]
:\eB[#U6AWW3UX()eRSMPJ#D+?T1:UME,>(X1EQ9V#[8OePU++aW;#-BBGA8?&JN
W>(UNe>?7Ea7F1MCMIc:SUd)d0<H=e1Ie.7fWdXL]\PZGC-g@1P2&O76#Z_)(@D0
83T_^eV4)3ZL:3D4+g[c[/LIELG]dK>bT1KSg3A;HBCX3J.&=GC1)]YN]I0bHGB/
YEFe_6^2J;:9&@g-MP?+D;NI+P3a^.9=^>.VR.MgKDL.7SI0ZCcTCX>)de5c37Z[
DcfRS?J[FQAdT#(U2]3f&K9eN#0^0d8,C.3g04V,LGG7VOJXP-YI)gX5IDESe@K&
92/58+/SBN9J3=0T9L(Xa^f>OM;LW;g3&_C_9PR,b<9OaA&&HW+G)A5Z67aLJ9XR
[e2VZ2?&I=UbH.DTHb1/Z#1@8T.e;2&g61I+LRCUQ;6&]B7==cN][[>cDDATE2V\
X/d3&@B4Sac.]4<J\(@ZMKYONW>D.;LQ<\aOH_)Q)XE2/<=c,a4/WS>^9HZ5d&BN
2E/I=B3[0AP9b6H=1@:G)W_K)#-eF=D21467\NcP7&ef.gED.eR6?@(ZA#TX7SC1
#L\?BS>/-P@dN:S@07[P]Z5DY8JC09&dC8FWU9JP-(AR.0ga[aCa_AZ=e\LE)-e9
#MHS?/GKS/@>W:;3R7&OgdM=\Ubf?7L;UXY26PH61KN.,.(PR\ATONgQ7ZBALIdB
Ub19+La4e1>f9-6-A:(M:e9W)WeT@.S;?eG&7SK]a?Z5aVdeJ23eXG;<>JMIaSKZ
(eG2W0=B,M-??XXG9KZc?TMSY5dWg&QKg)01c#5-RGZaMD/QY<X@3F8_Aae3WeVM
&OH+=e9ZI/@a4T9.BA&0BF1?ZFNAQK7QLe5CUU2g]/74accAeZHTGTgc\--gd^Ff
MP)7cK3>&JJ?8=P-M/[ca-7R6<7Mb+OG4e[K>#/fONeYKD<b#<1cS+R=<JQKEQ5(
<#.;5+TFC5bONLYf](:dR0Ze1bZ3b^YHS(B#)be---JDK,a9>ag3\Ie6X&a3U?5&
PN1ZZ[b[(K?YdW)>EK_?FZBRYC>ALKNKXa@4-M.EV7X75-N8d6VI<3g/Rc/3[;a/
A=]5,@bg;,dJ+UJccdf=dUWO#47;BFb(/JCA.1GFEO-fY^60FgI7<g)/Z<bYS>0#
#0W+X11AOQY.-DJeD8>1Ac^2^O-^YCGcHOG1L=6ROe;1T=LFS(;+Ka=T=+>PBcA8
4\.@==RT.)ORZ[ZU2)MgQAHE\aa#8-@CeBd\:6OQRE[O=8J#Ea)2ZL0)+;e)<B<;
<4gd)[]3GR>A;?2^(?SJg(@HI(\=;3X-b8&AKaJ5Y<6KA7R.BN;E+I6BJfQ81)Ha
_b)F/[WTdI\O<CR8GK:G78SVg2G2-[g<ZHC8(^7+;6.K8f\LR/,<e^U/-_cL?f\e
]V_@(K#B@B]7U[D/9<[LD>L7[=\M-#+JZObUH#Q6_F/BQZdJ]BP]J[/EO66T.GWU
7G:O.V#=K<[M5[0PN&1[[]E#@f[F+8<WGCG_YJe+VM.S+=TM=WT=&5U])D;&&/P\
GS/D1UT7<A14ZY)A8T^:d()9\Hb#BWA6Z^&(JV(S-BLIPWCA.]6JK8SH<;[&-#Xf
F\<(;d]5/T5GEC(A<_C#I#g3aK)PDUDV(aB2[d0LLRP<Y=5fbAUC),O(R0bc0T<@
/Tb,;0N<;//B555&DGgPL&Y&#&UaRL[JS+F6^VEFCdd]V;d;S&2@LX9TRN,aDcM4
HJ(^G:=O^)HY3TY,de+7N72Q_QVbWQ9KG=B>,UI.YPKS7ZHaNM+^.:F<KQg>J;);
8-FBSJ,^2D+?RBASc+]\^VSGWYUO7:dg^S=aJIZ?]DWY8CY15RCW>UX&0Ob&T[6W
7QK\]I>-3_DH=]E>T&[_?@XV8[CU8?g<V+T?13ZQOAN(X#61K@g)^Za:e.1H;;RN
C7O=dQe[d)\7Y5RC0fN]8EZ)H2]X3[6[GP0:\20.X,BT/^2O_5B(=SEK605X_[,1
8I>;OKQCVEHaV6>9[92VGbEX.9.3^:^MYdaJ<>].[SZa3.3<O^,ba]C]a8c.WaM<
ZIY>.:a1(T8HL1g->dY,8@MH7=W-=R,&K8,X\QE?21f+,4bTD.-FM#5-55@#U7]_
/E>+N&56(;VJJV<SLBc4YEebO.[M+4]?+YC^>TG^[6L7SgO7Z5.dWRKa]?Z)>(]1
HM2F6E-E^;Xf7P:F>YY-geIGD,S[Cd2-K1aDU?]Cd=E29K-6aM(QU[@R#UcGX05@
8JJF.+7I83^[(RNReQ1I_?.2?a;a0_+.4/[aUUBVJ&a6O.(^OHG4SA.W<Ef8gUW=
De/g[0O@Wgd)=^GZ&Ib:F5&^H4>T.?f<gU99.5bTdWa6@;6b@6(VK0-9F=OO8M@]
]NN3@0e^[M3HO[bJ4eN@I3KJ\[HTF3V&74TDLX_IULMYGCD?H0eTK]&OFY\3/_3I
a<HOe,@OZ-@X^XGa_3:1b(23U19TPH#1A3_];QZOF4+da/P0;4g#V=Z#W40+;Fg@
WS5]XSCR,(CSKO/QJYW7CeRQY,96DQL[-)?N_.TVV#W>dS7_.a0B^=0/Y=;P0R97
gDK?VLGCUf]:GU9),gIJ<)PAKMP^B+;;LS[#bOgRG_ZINULQJa[VD#PK98[gc@_c
Q3U]5dgOfc8gbP:--YG/\;-UK]YJ<N4<28aYbXH\YB:NET7BJfKTP3b08Q>bNXbP
A3e).G<&LJ>@-#L,&g>&]+V^T-GA^E4J:APe[g@44Id35VWZUOH2eR9Jg8<I@8f;
-dB2ZI6+0]\EU64H]/;J<2>JX+aHMeT36dMLG],MAK[.P??0ILY64-,@3Se#b3GM
a@gGb2JM]G_DIT2@Y>a4><CHK]GPJb@^VTQ)1BT8FGg<FV<Z&:fPA^(I::ReSe2J
H5_822)_H@aF/XI4c\AJ:D,)b_AM.M97XS6GSBbgWdK:#&[#+8,#E&ZY#1=O[V@&
]&IWaV1BJ1VA0,/@ZSW\X_e=]N=N;>I>DTMO1UgLIF]Dg)\g@0gee?Jga@5..I;K
>?12A7YN9_7DcCY;@)PUIe[H5/(686OS-J./>QEHUYW53AFUOS1Dc#CKb0;?gXa^
3-HcZ,U48[[Q<+e7^^HC.7>,Sc^>SgSN92=D(<Qf76I-bC[C[g[KQV5_f2\CdEOC
C&A8-8XbA+:(3;C3+CdXT&#U\e[RDV;Y<O89aEPM6-+ALIOHFgf@ad=@2?BWVYET
Udc,aUEe5f3LJGFB;-\(8fEZ,7@<1STG5@f2e4Id6BD>4_c7QSFZSF9BBQ&ECDWQ
9@D5aX4A6&JD3C6F\Ff6?g.#Wf?\F;</#S6bR65)\eECBIEGdVE&fBE4V#.D3++<
-VK+Z8F>Vg#4c+_F^VSD,P;NVD\>8TGfF^ecO0fSV;.C>(7V;6XP,=P^=J<4PZRT
^IY);\Q@CNaZd2=&<=OMJ55CC]EIMK2Kd:/V))_d5SgAH;VWFO,_S1O34973Wa&B
&SCg1O<&(:c,WD+/c:B87.0K\.E7]B7aLCJW)-<HaFf#geT?ZNJ7UPb<FUeH\VK-
7-F?c92&C^BS4(bOb[e/@g;6W(<PXXX(3ECHOZW/B@F.=J0C7C/PNeZO@V&3MH8F
d-D=-XK.6Vg:5F9)U.P:H0dbR+5[W?RUbKFJ1JH/aUP3(a)B]&0FVeK891&2K^):
G-UbQ_Z9fUd3AgfLS6SHOf7Z?BW/\7(M<9Y[FRQaTZ>9AG-9cF3]YH3R:@3OaX:R
@XOJNfDC2TM-,ZGE#&=U;RVJ+[RBP-7E64)IEfQJ#Y93=RQfd/?];2-.6O]=28JI
?RYO_9f1QI=X8@;bF27b:)[<L+<P:6<&&PS?L.K]8F[)7cN_C-b7(^<)W_L^(I[+
3HDdX+.@@_N+9K)e@>fN\0^7afe5+g8V,;K1DVFH-5fC@DJA)_Ge]KARLY+d;=LE
S&V4V+5TCB\C\GC2SD:)?6TADKeeW/1\8LBVg8CGWJ5_f5ODW16ZWWUIf6<_e07,
@2,JMJdbK9.3<e5]IX/^A#+U5Mc0d(dgcFF+A4J+BAN6=W13X,TRK#[<ZH[(;T@,
(def]_Mc9NWQLQRVcKD_QgUC0Y^Id-cbP-(A3]f\(ISaC6@T]PE]BLI0&^_NeM1a
M=#X]VU[WA8a:7<bM&-ON[363VPEAYa]Z=bgGa6:G#@N>bA.PZRQV=dD8UEG0NAf
GaD&6Z-)ZHRP-=(7IdbXVW41K7/=,QP].fUDG5a,(&aD8a&7:O^c5]VZ+,=1A(R:
1?1@Cg[UT(.MX>9IYe_@L;3\8=LBdZ,T\fb8[&Ba^1<[#G)g6c[b0E26[I+]aDC1
^L/Vc?T^\(..=UgfD[TKHF3DC?X^bOH_,@CK<HSAf7)T5EK9S@7IIO0.^;;<SW^g
65N-SZB/WV9SBF\OQQ<NA2Md-GG:+7T&cADa3+,\=PEF2]FY[H_#=1_:a-Be/E0Z
^06@,A1\C<@MKO@5J33N7FX&0A[?,c5SW)6HK]Ube8^<CF;K21([AJ;gJG9AKL98
KM,.fE)6T0Q>EOQTEMK>;_(.3+W;V468E9C9^G/TR?>@M\S1_+Vg:-NO/5+b8;?>
FL<P&CKZP[U-AQGf@^NM43_GFMIV9+M0MOR^OPb_6=TXZPT[MfV^<)\6,J.+RZa@
KW(+>Qg;(N1UCW^<0fGe5c=[+G.H4e1Cf?S\23_d)1I[^LU1CKI(<Z_8.cSbGGC3
/035E.PP(<7Od(O.C<4Of;Pd[.OS@HNM2e4E#^)f?N;=fN77D,\JM&;;TdO80[9[
3=H[H\:dV@SEUUS_R#L7^AT[ZQAYbI1L]\??P9-N\<_cbZb_Z^S.X[>ePbe7c25S
<DE@WI-M;)I0)5Ffa(H28ON^4+SPB8<dSD<(UFK/?]64If;BHb(649Qf4P;1cC-.
-fd1fYf+UJJEJGM8>^+ZQ/M\7aRJg1<,DXgfab?HK3XDFA+4dCL^>G7,TRf^K6VC
/^5c3EQ0KUR&e7)109dEgC;OU+5E(^Hb<N,a^9XCg<8FFa0VX:D_cWV-CQ/NXN[G
d,2a)&BN]4KHY=+Cd3QZTGB1b0[Nf-2Y0d7ZYIeJ4#,-?#(I-L<+R35aT(AX5\?I
BB.ZUQ#F-+JWK=G[-3,;F(@gM-WKb,@P\)FHFLc^Qf-/XJOd<fM7(<O&RH78/Z(g
G3W[eZ-5M<1G\,XZ,_-1IfOCLR7/56PEWF&eaV/1+,W?H:cSMN,ZbWfgCO)=R_af
QP2JKS6:CF-JeY2d/:;A3FTEAf)EH5HL0(>ZgMRSa?UY73B>(+VgB/BgbN>V>H7Z
7e^,bH5YH@X17<-L^MBc]&LJR]ad<ac@Of:7^AT@2/)#T].,KZ&#W7>8XM#SO+XM
#5K^M3ZE]7bC1,]G7(SG\CV<S^BbW>f]GY)X]J.TbP-&\c2O[+cE;HN.M_Z&/ZFY
67f]Yb2:Ue@^W=>=[TC/Fg2Q/Z/\2DZZQTE:S#gG]CX@SR1P\R&P.a+W[FC)?X?5
GW&dV:8c3_V512G?>O-dO3FOOYULW9<M:H+3IMY5J<e4(+>21VM#fJX#M45\-?+c
ZUa-d2&e/cD^d5<a;AA1S4bH,=E8,U4DVG7Q]D7)_L:<@EHK[]K5T<e-:<N4B8FO
E:X9L50X@X+1E;Td=415ea\Y?NQ]>ea.)_U8R8b7c72OB)=RWL^XEe@9WM<;b#LW
LGRaVN+1HO]WR-^39>8-52=(S:#H?BKAE]EFH)39c?ddXIO<>\P@fC_;Sg;G2OYM
X;K^1GbZEe2@gAG;?DcWN8O;J9UU8-0^eM#AcH\McNPaZWdG1OIZ8]8.Q4AM1,F=
C;2GR_YgQM^ad_KF::TQ4fBZUNO#>8[=\Mg\<K]2bZXNM^CA2::=LAZQ^W:b.R.^
D6(-;e:).M<@&YJ?[RG)f#WD&bbLO-gN+V,)30b@]1W/2b.1&ZUE[K,/,g3J?b:Y
g9V=a&FXeV1OX-)3d7@3+R35-<Ze]b86>T(&+6<<cDZa^O4CPG7,)RO[,\^V6MA/
3X[R=2^8:6NW]]OXL2TZPcJJYA1WQbW(7=RROg7L\;+^;QIR(5_Ig^_.&:4BOGK@
a<TgE81JU>=&52V;<1Pa<c)&GV:BSP=3<^WN/VP-(HcNeQLJ#);(SB=)U[CET-81
Q&V<7E&#bOVVYeS@N^(Id\_.FQ7FNS=/&.,WHC;3Y+(C5M,#cVg:@UF81[R/9Mc:
K\[b]8T<Y7C)2^(#+LW4C2cB06[,gcFg-#P3e/Y_0@)6H\7Q.S8PNK(,KdPO^T_1
@K(Jc07TL;c),/[&5N3M+\bI.8:1>/K_\+PN9/HeUFPR\T+G^J<PC6^\^TIec/F7
HT29T:K_V[Lc9&aNM.IE;8E=9a&W^JEPIR<ebG=1&B&6O#YL9&0?N;=KHA3[C/g)
S)BOb>5[OB#XTS#<P^CT;JK]CYScPc<UTG;>fHdcI:_V5.Ff?b0>/DMP\fA#ZfbY
;cFU)MUI9-BG^UWD3XTeWeTBIBBK5P28H]RcZ,2M3ScK?(:bB-=TbJV3&g0P[1\3
_LX6N2\BFYe_/cA3)^XT]9J8VM<OGeBNMeZ@b+4IFUgVP_IBgCK[&@5\M]KZa+R_
4]#)V[G3Q=eO/H+(RMP5VUY+C0Q)#FH8fW^Wa=NEgI/H=P<>/GfM<^3RI8BL^4+b
2<->\T7V4&<]_]IKKDYSXRBaS?8]a\89g(^15)\-fdf+7B,.+DAM8[WWUa5cf6_X
[](N^0)N]#b+9^g0[2O\QW1KHT3U&7.V:P(T<D@f;9/Q9_=fY9UEJTd)5I#0YYFC
d_MY_CMXSY9GBGI4V;d0/U/(7M+@a16gA-?4II6_O=ZUDKNPQa@P.M(X[V&fL?24
2a5B3PRY]fW9]74IeTeBMET5RS+P0c-,8>L[Nce-G3d/A^g5SLL#+QZ\3.VZ4-YW
(BR2ZE#SeLWSF6-1G)H=]@TNRWNC_YXI\3QTe/GI.I(c1_bUQ(d7,e?>=-Zd=f50
MgQ)^W\3;Q_-#2+I)=PG\\7EH/A/0,#V5J</HV,#ffW_+aD)(4bBXGDC<[XD\K::
B\07gY^UbO.S4LfI1R9d,/L;^g:[a(#4HPQOE-3=3=B^O2<Aa#SBN<Y4/_192Q,c
XNFf^J8@X&^FSAg.S]=WcL7V&2?)J,;<OSD]a:05BL02J5Z]M<O(^LIFAeK54+5V
@Z?P3OFNGTEL[HC_aL#gYWYI\;C;Ee9Qb]cB6&S0,?XLe+GgJD28RLMTZI_,YDJ^
&MKB2&Pf7+d&VK(_J\cH2b(VdIE_+9RPB[IFaD9F:K&V1OXFe\:c6G=FH;]G_;^I
B<9e(a=1U\eV)S6,,_R2MQDDa6D)Jc7-4_L_85AX33RX(.LHMA>ePadBO,OEL52,
GJ8ORR(O.YdU4W02N/e7,6K+g(be;(eA;4YYV4NWPG[J9;)1YgIYQ1SUU?<TD,#b
M041S\-]f5[2V29FO&T/FNLO1=M@be5HcC;gOD/dXEa1]2?+T]>+ObL^P06a>De_
0VUV]LOR31H+/ZQfS2^D-+1YaF/3&U_]ZUB<\EC#K.Q6_3d<O,BTaLa/?4\26XLL
A4-D#CWX<=5HIGY0f?R#B_-4-a)V6N3fbQ6N#(T.(8cUKNF5Hf5]U]G:N\7bN7Bd
,/L_E6CGf4R@U[(3S.ER?I2Gd.O7S6;IN:cf6,B0U^UF?)6+G[R<PN0dQK6/42X<
ZK]Y)_SBJL-XIcC+1VeRY;7-dZ\.SH.K8\&@=;TW<0N>YHa8,gL\Y1BV,b=K=S[7
3C?Y>bHOH-/P]DI.C5,HLf<]HD95ELHH1,YYPfV]U/\3)N;af1Ic?Y@A\^,/5R=E
^DMYB(F9Q>3IQV=bOVBEZ82DH(MfH5fS:GW[_.HR723I)V39VVFcF=)]5GA6BIED
CG:.TPRb7JGB[#1G@fN4>(8.=4Xe^X:Nd7/>N,)S_#I@Cb&]^E7VC7[faUMO6gAg
N\E4J\ZSB?gEg)_Z]cVCX^/#dC-#W<I@Cg:255YDR\FUI<KU2f=?#=#MIKH\.=d^
C743?.ZV#E^&:#-;DGM-f/@.B>If(N7RTO?E<:<323;106+=/&cW^2I(44Z4TW)e
[;OGL;8X>]9N#@X0d4D:+?;:S/.f&EgBL&&gFRI50_W\1Ue<K+[:+e#STQYQ+88#
XPTO(J,LI8c^@e14cEc:G?)6=(O=FYaTIRX3B=dg>18b/WIfDAH),EgeHK[3H(<3
O@6>0SQ+af(26FBBJ+SSF2dOC0Z##ZfUKCU/#T;1@+:L4BO6;?DJEHLO0W2g(OA>
4bV7M(LEOZ]e;B6VKgY#PQBB:c:-QbFOd<4(9G,^IWg3dK/L2&-F^&a365G=HW_3
#YG4(a]L[[S_/N#b;A0C_4AOG/@UVH5&M_bf?B,W37?-Tf7[M6CaKO\WG1Fg?0cb
3B4&E0GN.B.ER0AWMc)7,HF;I(ZEZS5e-=:^3XB0<HK&<WR#@>RQ2+dc&f@5.3U/
bD.E.bI8)JU4\S1#NgL475_V.2HV]bLdWYBXaEGHN57OPJYB)VN6EYI6;DNG64dZ
ObBb0>R;EIP:E@@_]a+@dDXd3c:31_4YF>]IbNFO+Z/Eb?.#Ra#8ZEV2ZZU[9=gg
fD;ZRJa&aNT-g?3_Ua3K)G5-;+^KaZ:37#IfMK/PF,c/B:db9eHR9GA&_)RK(LM]
g;&BVcVe3:C3:;24N)0;K4Y_J,eEd]FJIEZZZYg(9db5D9D43ZM:1/>_R14-9\7]
TH_4D.a3b+XY1#E[3KUGN.2A9#6GU+#8-GU:^Q\Q[DaQ;7IO[VLRFDAfTb0JMLM.
3E3W,G5?;#YZ5fPSN2N9+@c)87F9(BI_?G,7/#=1VW<gHAf8544<&0^)9P.c:+M_
]BLGRHY)U]-,[S&V5;/7/+\DP[:ZTJ3)7H3GWJ^]&>VFC/[28[=b.0g?Ef[[@E#&
79g2C),M4Q;O]VU:=e+HD1L93/:0aZZ/fW]&eGH0_RK/eX_#XFb[:_5LF+JG-Z1R
,66bP5?HH9+D9c3_O<2S8HcIX.UNBR;S3#F.;VI&g^@LV@fcP4MKcBO)Z2ZGC:MY
,8[:g+B@@H)4R@MUW)[Y.O,OGT9EAKW;/.FbF=>JK>&YL)dGe&466B.R,?0[e&gW
CJ>@e2VTHK3aa-\[5045>-P(^b;I_QRdF_N^\JT?K.YJX6g+eR=4W.[fS8+T0_(#
>A147VUC<LQKW.>5FIV7?2NQ<IDbbfL>1O0PENfZC<Ed&:3]6dO3T574_979,-43
0.c/PKLI]?8a@TWKL4cI:fbDWAfJ#aa,7a2KOMcY/,H\&3=[H9HXd^c61HQ;e[LQ
Zb<?FeBQ1E95PYfMA>6S+=53W#M/+2@1@FF+)dTG)Q,S.O2@:+a[6_<(&Yc2VAU[
STU+MH/-R>Y1BV-J_<@-HAN3L#;D+c[bdJK9#;S\]\I.-UC>4W_G(,Kg6f,?L=:(
LKNHe0VLYKFf7U3#5TO+7SR2)MbD;=b-GEBE\(+H=,QSS6F<;24eXO1<M+?@2g#7
eYJ#]MP(3+<.d+^gbFL^3O);[T.P9adAE^MYLK+4FSULGY6aeHOO<O<(8GV@aVG:
#6Jg/E5;T#D?2>FGG3L.M#fK08Sg=7?62O/eS#=R0YV75:[5HX_&f3MFOVeJeQ,\
T#VA7K3^KI7.[GA/Gf^D?Ec<M2aRa4KUV:&cVRg96?FH0ZK(MIP:;C4B>c?b_F,/
]eD@&;-;L3ADV1565NH3?//+cU9N:=9Md\TR(/P34T&SB&-:>Cd.S^/f2[9V23D@
99ZUd_dGLaSefEXYO&A&38;Cb0;)f]DS3ZG^B83CLX3P/1[)@M/LT16V,(@&BO.U
1#,CL.:11/0Z+TS.]gH9XUd]ZG^3dJGIOe>F1bHGRID0_>c\M:&>DJ8N/b]-TD,M
T681R^^?V@XLg(7Pg2TEeK5FTTB2VQ?I:+5@S-MP,Y@LAREWNX-G\VEUUe8E7ULR
aFDBfGA4Pe4QKYNX7dF&:)^GCT33[JWTbB:VTPdT@(PI;I01RH^BbX]Z\8>TC_C3
::4,JTeDcIbP/RR,fK[__&RE>=b1[I>8=.BW[a&;OJ.ADdHXNF?+U8QVTT2.3YPP
U[L-dT@a0\LU9K6MW4B?L8->U];^NRS;C\H^A-9<)=BeT==+9TQA^8;P[WJ[cL1J
VSH&\b6H:[V=^=YMd9N8PbXR\IY@OH,WVc70>&-&)ge]e:d93W#VADJ\#14:@N9V
_G7F6X?<af0FgKa][baWbcG/@)AcfX>+3f@AA2O^EM?4Id4YU6QAH)/>[G/,QT+/
:2+NT3d2I[1c=cb.;5X(AXC.HX7C5U#D/fFIgcWZW+LNQ\Ha(aW39)QO_PU?/CXF
F:(>[ANT#33Y1D,d1dR-&(D^?AI58b+N>c3:+4M,&<]R]EKUJ]7T0eQ1B?d@(afe
d__cF0V0YF=^8][[B0V)4Fc^a<Q3WFF,Hb\17^fE5cNcJa-+#Lf@3R9&/Wc)<;.7
fc_a,68deN2R,4<7/U#TF^,dCR1e?H[8MH,-B;U8c/,(J,6(U;3XK9]FP4HJ(aXX
b@3\;+7SU\(@P/f#B)^BXb?GFUOg],==TW>.OeW4^9/8)3_bVL=BQ;?@Rfe+:,#D
H7H+5\(@BcX4VXeAf]39>8,6gJ9?3,<7K[Q\KSeZCTE[A3>91c&5&N6ZEZ@\,-b?
3_,LQRJK7T=gM,1f,8KcD/RFI-W5R,ba15IaT@STb>/Q2E764=MEB1[&^R<RT9VT
8L@>WRRT7N^]<6g/#2WNV+&5F]1)O<^4I5g]b/9K[d)N;P=:H)1gZ-T5X:Z,fVWX
PSLO,+=^38?O3ZDP?V5X1VdRFF7E18KU>d,(DXL_Da&]a3ZB05=gQ_2J6F#_bV(Y
SL4d\=+.\DcV\]9gaD5F@0?E/g/^RUMZ&5gR@K:RbBZT[bU(cEKfeTT6D-_3;LT#
4Q;M6R^UG9[Z;g[XY.?(?\G,FTg]+C,-B987;c8<7)2Z8;LcQ44[N3F)>@#YA95:
U@aZN2Z-?6A_dd^_?#5(#c=ZXe=FAAbJgfPgUB+)e^PcP?)MVE\cL65V?D6#A6bO
cg5Q6QCI6M0;g?PZFPWaRG[bc6Yg^J>,)+c@7HJGe<a(aXC2a7[>(\RVR4&d/dI,
5@.P3MDUGBMeH-UV=[QY>PDW;(??TWTM0+LVKcKO[/DP6(0;.4OK<YfKHXSGaWL#
_I)af0=3?GH:aR+e)_JWf;557a;b:VDZR+6FSSDQ9TEC8^/MM[@MfGYP\VMTX]KJ
0AF1K5FZ[8A-E[QbB:4[XELP^T:4E]-,\GEM<K]VJ;==1F@ec3[Fe),MO>)LbOF,
^,Y&^>:g#FSI2Oc[@0)0R_fFdUS[Q;Q6=\GQ(6(Me\Td4UKID(2V9KARX1LLKa(f
G8#B)Zcd4g)(?0c&V18cdU&4&8B2cU8(g#Y-UY-YV+-ZKWU^L2U53\SNX/(:B>W6
b,g=M#3PZeA,&_Pe?TGU+IUV_?Z=]=?DdPZWNc6R[E\6F5AAUg\HJ>>9RYR/[F\@
eM4H4:f&bJ[:PM<A?F5\d89_2J=Ma)/2-](LPNCM6_\X1BW>>/\V;Y&5gDb;g=dd
&8,]+]LA6U<1YFE#:e_B3V/d\GHaR4AS2YFKf:H5)B,G3[](^XF:f+7e/5V51(^Q
]EKTD(K?&Q)BAd6N-^ALLK9C0Y#HgWS6.&<)VX/Hc-Xf6F0-=WSfc4#C,+)J.B^/
NAaE#:\#):g(]^/a+S0X]Q)S]#Kaf<K:UH7+,-QNS,FN:)RDOAG[[aRbF,DJR/5H
/4dJ3M:a-R^LF0c[ABIREaAI.ZVV9b8)H]8ZUN?If3IK&C?/A5I#)#E#.L3WV-b,
I0TYA&9SRT,SXT@a#M@0+X?DX7&NI#W6CSOgU2-1MH,95VRSaIQ]7R28[,1Q+-<-
MMQDCQ+XIMe]VJd#@bSQ)Be>S&\9>RI0@fWCV(Q-\#?R)4bE&BD&SAV=,C:NW4QE
aJc;IGNSS,Q)SM?XGTN1gY>DMXd97+WH-g+JW6Q2VGIKL>D<e6=<dJGgA[+]]@gE
Z->R3FHI5E7\1Oe1QG/e]/CgD)4.O<;5W+YHCFJdd&<-O92)e7&;<g:34NUGZHGX
?[^LP/B](N;f)37U9YS;]0Q6cg+gd-a63Red[_LNQLC8T7+:E3UPNXFeGD6649f&
aXeWN@C(BMae5OM/Keb:TY8d<0Rb?9KJ^Z6NMBN_WXA8#M];cPG^,I#(</#;bWFO
LbgUY;GJW=\c?K(+Zf71S7?-;#B>42O^7[SeSKd(O:aGTTDMI(AJ(UR^4(LHd3<T
K,8,W1[9=.@a[8be@^\a;QYCOB5AU&W4&-G^=W@JQ?MINC5Z79XRafEA>1QBSXV:
NR5FCIANST>KD/73VZSZTI&P)7\+]K.F.1M\CR_dD2-+XJ38L>DSS,gF]7M6KTP[
8H,.a@QF//U&>C6@,#2CG./BeX#VEcA@d8;aJ(5?NWS43GeFRWZHg_)>8C-33#=E
JZH]GE,<b^;g3Ze.M\@_3@#2fF#]UH563@bF^L[G1RZO&3?ZIZ71Xg4VA(N3PB5R
P/+#\G,@C@VgX+LF^MV1baa2V=Q[BPHTJ8/+]^cMHEN>6^UNX/:e8VQ0AU]S5(,.
Ud64@KUSF30Q:<([Z(XGe[=>LOaKR.=,e7NBEG)MT0e:SRD)GUdN(R78?;-L9;)W
SG(2W38O[;K8B8MEYDC8;YeUC5b@:,b8>FG848S/:7W4VNG8GHA:58@dLTgI[fSR
Y6GbTf./[IO<.P^D(_U@+SWL\GDL_IDEc@K=+I?SQB;10I+I_1H3J+OgG#V;Oa3K
5WPSc=X.YDA+XaT5?d(EgY3(2X.Mb8H>KDg>bGOMZJM&&cU:b7E6;ITaRe&Q2Za-
2T\,b\,e?^22B5_L^3XBVKbC_4+(>B_Q9FT^/)aVZ_NCGb.#+R>B3E]\2?\9a7F+
>;TFCGe7M:f-1S,CI)-^-]C_M#YQ0>#,H+MY2AWV,K,ZE#(2:Q\(Ag&d&NWNG[/5
O@?EGU(aRdQA/CbE>++g4DeT8fg^[Lc@)C@U7\IERS#V0LBKVI.P9HId=X519Y[4
]bI>1K5+eX]5:f-I7I5Q<3^+Y+Ja)VM(FNQ0MEf5V_EKD==bcX2PG8\;P^0JI^&K
&2\ULCG3V;:CbegFbcI1COEGfHOe(E<B3E9L_D3g)?5gRSC5Z_Q93_]-TF]Z7df^
BF?54dS4W^(bU]bKdb>T[AJ8(X5Xa,QYVG#7Fc)^P8Q)+\L\;4@g(a[\CF+_0I00
=CKS^A2+R-Z(/]OJ^[4cS:I62L6gR59;B?QO.JL1U@S\<=.)F);d/>HT)FJ@_Xd>
LfRaaCSBYQQ1ST&(E#FR[PK,ZJT@LgT:\)Sf^/2F[(V>;OZ94KXU5>Aad]3<N.dE
YTVV5&(bLRaR(])8fFM<OQM2baWFVJ0?#V&,A8QSd8TS/7DCY=<&f,K+WUGO@Ca;
XLbHCF2F.LA1>Mb\VL/)3XWU;)>V?T(P\LWMc-B(<6M1ddYWC(a^&c#:)(GWVe&Q
KI&SU&3S]/ePRcKROeb/0.g]Q50HT@Y?PfPS]gRe]R?(&+Oe_f+XJ&^DM[F(,0NE
^1.=[/&;@=cW&E1b:4RJ-KY=4[09LTUId\C3TA:fP]Rb[49\]E?:CY>&Ff;df]2S
Hda[?8gBV5D5dT-4.7W^1>LG/FHPU9(:@#ddKdH]?V<?+@=3Leg(,Aee3NFU52S;
_V0.>(5JFgPKD=b/aDc4fHWJMG:88,(/?;g&YH09HD-M5;f3KY,a)381SI_RX.2)
#,:S_Y-9:T#43#.)AT^J56=HePaSU:54R=,/<^Pb9-T:?c)?HPQT/<XFX&)ENcYC
6,9WO/=TSQ>FL<@;.1E,)XSSgM.7_8bYXJIf\_b@e5d6cL&Mf.1@S^M9(+)dF>T0
dWFfJ(X/1\aRa:TX24DCd-c\<)1?MHC>5ZfXH,UA)STQTZ(.(0,AZ)@B;;AU:P@N
Df@&W<Ze.b0dJIJSeV2<X&PId541X]LQ(K@&SNS)TR0RccCI5,O/55_YR7aW6SS;
f.5U,dJTTa^H\c,RAERS6)e]BdgUVW3[6XMB8=X=f<U:D8GG[C9:?Q2FT4)77Fd>
&DC5A+7B(5JL47GdO.+\dZe7<E.=ZLGE]0LgI58[89-C7)L,1E^H00^MM[WF-FMA
+0FeHN)KHMQ(084YU2Z31W2@N8CS-34C_Mf0HbI1H=2G+F128;1SY,GX>Z-f^NR;
6W2Q\bYCU[>^+c^6SDI,,G1W<B&2LD4):4-Z.[g(=f,d[Jga.a1a+fEOcZ,?gHZR
a.3D9RC1C,(^N+[O9VQ/[B,UR0(c)(_OOQC:T.5.8YPFE#&);O6,0))+eb7V[2>P
J2W-1)FRF@OQH>f5Ga5W3Me0(5OYJLQB#,N.ND0dQ&F;T<c7L+AaR07/A&53UbeL
aGgFR9-T.)5,bYWB^b:ZV_d)VJ877G3gN]XDbg)O-++;M?TUCPY)HdXYL(X+/5K[
V2;#JbXO)1TV]74__/3TP9.K-#W39YW?XHSBHa\<FYB3@ZX3Dd<?9cCa7TR5_K)Q
V?eg-c@G?JH_cBC.cGVV.\J4\Y6\#\X4<S_b[COKF+?32#^9@_M2QdATdO?bL4VW
VWB]?G?eI^E7,b&RJ&479<K83SPJ#K(2(Kacc>&1fG_LQ8DLX()5O=@cF-8#Ia&^
&##6\6,;9Aa]4NV?e@MgH_4N0g70d#9&:[;0S\\D1L6TN_]#QS@Y2J?<)=7>5?RS
PLIA^76>bI1XG4SUYKTMICg;E5->5d)]D?S94XU]Vg&YY4WNO5-A/-/^(<M(F:/<
&^WB:A&5N3W)HQBALKE0E7.2CZHF;7B4d>\/CZQ_/X0G8KO7TDb7)M8fF??PE2M2
\X?gEKHSc,S)g;X\<1@1G7RW/?.<:4f0b@B99W8DHN<?Aa3/[Q?IebW6)De9:]M2
WRMX>>X0-M:Ne^.e.OEBcFb<_V.2MgB42-HU7H8\b2+<09FS(T,T\[62AVJ^KaFU
O6,eB==&@3HL=5gURY[A1PW+F,b)4HZMd)BQ>#BA<KC(Q9X>@.F;-d\B(/8NL35?
Q5_,#HJ\\.O&\6N-@gYP-9dSHHP^KB]M#PYAabCNZ-/>e5I3Q7BB^Q#>(;a_E^7U
21.FKZ4=K3T?08LUWL\KR1P]Y?3(V])BaC_#H1dMWLM#T#]PZ\HV+a]9_SLOK_+A
IY475EOa;2fCL\EP3JUSJJ]AI^XH9Z^S\RB@OFCGAfEL<]W^aC,/YJH8P/E^9B.L
DJ.IH72,N+#/1W12Z&HeB#\K@LfgXd.FEf_^_W9:J4@GfT/<[C9b>A1[Q/DaV8>B
)N.L.Jc)d4g-+GC[#g&XU\C5.@?:.TA/5dc.;-04+#g006?d=K6_+BD#E0Z<>G@9
T79_2J3/?)+a#6Pb#KdU;5(GS2A978\911U]VK<GBKg]98:Qd.W\bd2-0U;M>^NL
LU]0Z_.g&:8)_8YDIU.SO&Ef)H^Z?W3I\V=S@15D..KG\DRdO?T=eRWQf<aJ_9)Z
b&Bd<F;[-fME,[_5LSc@0&.)NDUPNJ[(Sb3MH3I-+-7cUNO7JeaP9Z[N07IEA3b#
eE5I6?+bFdCONL(BXOB,./ONWV,7KXWUB28@WJTSNG(GPTWFJFN9ZM_a;#2(#IYg
EK:d(0+M;4+g^QeD1>0?HeEG\KN:LJB</71JLCMUH?5O9:JcF3G-d1OS/-B2^.F;
@Sg@TB1ON>X.9-D.P7G[UVDAFMJYEQeO)HeW#G(8>ETKW(#MP4e6,SDag+:>A3fI
>eD)O5^NSW-^9bUa@8_SEUJLBUR3[R,#Y-[X>8Z(^;Mea@HVO7[=9;C8UEa=P2ET
2KI&Q+,QHL:ZPFZW5)9\I89K@f^b4[ZM(SQ/OYM;LS?Va?O-:/_TF?ZUa0<#ZE/C
&:L)6;J\-^/d1&=X6OfH#C?A8R3O06#K.P]M/4,J/,6[C[.Aed7<B3M&5&UY]3I8
Z=:Ce(HCY(H,Z?S6Pa\.559V9KI8S.U:MKdPg8:1eL)Q&/?PJESYRC+HHN+;2;BP
<ZZ6Ib_O=Y<D/5H\KLI+gU=,TM]HQ\N]D9]+8\?V0SRCM0Tg<NB1T\]@F+NIY^Z=
,2Mg7V&H[U7M8T^]LDB=#)]Y99T4a#=Dc5Ve<b>E09adE4bURLNdW.]89\7E+K?=
U1(,_eNaY2ESP67:#L);&dKG8?Y7J)ZH-9D,G/S6DB;9,WFa/dH[7RO&/FEQ=@86
UVf34ZFY#OH9#W7_K0-(.9[AE]EbXa>A0@UI3WU8EV#a-]3Z,;L]9SJ=_SP0=PQ:
3#B4?K^5W]?GS]7@0<d7Y1AYM2T0c^&\[V__[.RJf:GX^Z]:QRT>dXYW[\>aQ_V+
<e,&M7.7[T,+eBe13>7HbDL4&VZ_GWcG/eBCTIgN18IVI_3+#IeR?6cfF5593\TD
SH[+/NdaHL(B//UF?gO:7Xa:,3,V.NdSE^RXP_U:KD_:>QJDDeUEQJO4W24:g[:7
f/&(8W[J@EKB7[+SXOfIIU.L[9#,KH;N>7AUUD61cdc5+V)5C.ZGf5;PcR_\R1E/
L;;A-WcgW+]c,R9SOL2^SY4#DX[gb\?S</UH]2HSXE^/_;I@1IaE-7NIMWEUQB<S
68L/B_^WSCLccSP>-+2V5#?/=U=J/a961-S^&.J[:W1dEQI,UA(c&1-Y_c;R>:W0
)074Le6b,;?6Ad96&,0K8I86Eb/:O&Y?a(#RPeaQSVI[?_>7ULI#7&8;0MX158AY
G=#A;?[;E.6fL+)dGEURJ56ABYVWC/.U@OZEO5&_(5M&DS-Y;]OOYcT-EaE]1Bcd
<Z,a6e/-a1AO7<dQFG0ADDS_H;=LUYXEH>OX]2[IEYeaN#.P88dR_[gD(MUa^(-9
7&,MP>2@RZDKN3(;F.IQ.@4ZUGW?QfXbGZ464LD?QSeW^HWG>;LJ2OB#,>Y(O5S2
E1>8_VP5e[Od3#[+\^[aWM4LfCVe[K1dD+?HNU)0B._,2<H_POdD/5EV,3:NFNde
d;W<K8V0(@d[O/8Z:@CJZJ=]5^_3QJ@WYDA=2Rc)&D.<ZNEGY\eE6C2dK8.XC&,Q
MY&\I+35:M?N/<.>K/+:fB51+,:?O>XL=K8:8,@]Fbc6H@U7b#++&:<#A0#gd;>B
WD:O_MZUaGCaK#)&RIQX:^CA0]dE_?]H&FFMfS?3:<X,KN4B-38;0-(1FOJ4Q30[
M<[ePNYX@.TKSPUOVGCFg:RKKX.)UM3NAR#(&E^(K\CD9NW6>@>D(_KSA:&dg<-:
C.8=7BF2GbO>A.6[;6c07C;5b#SYWa3^dX@EHAcOf^fEFaF+J:HHZLJ?#2LBLGRB
>)2\6Y3G[M(QI,0Q)L2AF3LZ4,<.M#LfRS+OMLa>.3Rf&TGBHX.DK?POMfXKBM)&
,=)aI]6U94R\+H@U_DSdU&6YTJ4DD8(9f53FW;NGD+4^8c]a[MFDcL6AA6(:I3<(
3.1I.L^)D.PE_;WPgH<C,U(OAIAII50A:F511.g&[09?FT?&8C]:b,Z\GPZ58AB;
H8IYCPAK2cQYISXRNCFdHUFAF>P;&_V=3H3H_g7e-F[Z5F?P3#^Z;&R)-:66D2bA
B?d5-NO,B(ZA^@N\ZLZ4)XX/0X6b[#H?O5=<I<U54b6G_?VQaVI]\Y9a_E)3LP#]
[?294BQ&]5;NBQ]c\GM_=EJGE,a1W@@e5,0IC=9YDK<USC,FY40V2SJ1&KDdQOG?
^dG9f/QJ;)SDXAYDL3^BYON[T5A.2Y_XV.c6EbC@\WDO4aMN8Z()+fP=AWTaKZEJ
IDO==_^=3ZL2K[1@U/1@&R)Q/1)\?TMNOPTMWg<I:^;0F900V^U8):B(:3^8@dNb
X,d4#G-I2B7<+e&PW?bLS5^e6R/-23&;E:##]UV>\G()COTf]F1c(1Q35e\@E)[T
3aD.P3B1Be/6?IN#C)#3W>@@b,])e:?@V?+/-&Ya_>TB8cQ-S=R11)JS6<FLVY#J
Sc5>b(^>.Sf:B0^U#@B9Q7YO&bb@<EB\bVa=<4&e/;/63>AQN(#8d>8;2GIfba0H
Y&c8.G(KO;5IPW/<8)7d69M=Y#B+MTeHa6;O&3EVZE2H7[M_@1]Xd=CLQbIg?/NP
8\NcJcQ_LPL+cKA)E9^;e<XT@Z:OF/DRW[\<^b?CF8IL2OW.29e&NNDCJ(5=/S0B
YF<]6.f^;5<d\TU:fL=LfXS2C_YT3.9G9-R^0#>N.68]3@@.FH@ZY(VC]Sf&+>BL
U\6(X3&VcE3VU52Ed97M3[ROW].cc5S/:a][=KJTKM#?)AcaWZ:^S]+S+S;_FQ(D
QZ-:M9+#[#.dMcU?XG)#d]QRL/MeJP#K>\1311/c83]93.NXg2aXO9SKM548#_FK
IP@X<43Q1fA3Z0HACS6Qcfa[d4GgR<5bQd7[/]2UD:1+L>6@2)>)^^O,@110&=YI
Za.<7QQ]>N203;890\Nf56DVE;9#Xb\95Z(BeTA^(B1R4OY5J?Qe21R0cV/^J;fV
DWZ4ODYK_;K&C[]NOC@H>1=I:AS5@8J_VE/1K=<_(WMSI<B^2TYT,=W_4/VM?]8B
-QP0d=NA0CC_NfIN@\-dZf\f6(e.2?.8)<IQYMD][@Hf70U+\:3UBLQ@fc[.,A),
RNT_+_fWG9=g\-[UC(<=WK[AKK.f^c\cgXP;#c+;Pa>:V^?[4E+\WCQS@cDX?1X_
M?KPT3++HfbBXc-M<&[a#=/QJIf&[G<f7RGV5[BcWM7f8R5R\RGZY>.I:N^KC?:,
GdBG0H4+=A>>BVV/e+MMP3KDc<Wg:8&9R^MHE76IYd8]</RM<3_++-6&MJ66PC7?
X3Qe=.YWTERTV5aD-^d9&LL?TJ;7C??TUb=g(M[MfVT?b/+MdKJ/fE<4QFARFO.W
9VUF7^_)8]SNOS>H8=51R3eHaVcd=7T<]:DN2GGU+U2,,-R.P__Y2Y@B/U])9>6;
LR^a&[A605@2=SD.8=YGSP/0:8b2H;gNK3,F6\#Q>dB5\/BMQ25W#RC6YWBN?eeQ
C5-D(P;@YYV&d/40dL;3,:FM?&E4TA>XX_[PVdQ^@&,H1E]af_<0cZ77a,N@+32e
UR@-_I-MS_bX\8dc+S4HM[529)Y7-gb[K@\ff>#C0Ufg1B8I1ae@<-=TRdP3^WfP
]VR1[cEUQbZZac0a2D#W5d@\)4(P=ES\VaHfLe9\cI,d)INIVS=dEL\7HF3T:N;T
MELV6485S<c7J#dbL>]GA49,G;D#7Mc^_eCD/&F[,QL[G6MgX>RC?&aId4KV^8+Y
Q?/IU=/W&QR[&(YaSK@[5.g\9R(/=?B_9?2^-eJA+LbPVY)5V4RV)e,.2bPUcT;0
W<M3<C9OD:?[X^J3aHAXP>OEdPZBAObPBU;Ka9bL,)IIU:6^XDR;He)CG]OO(V.(
25ga8:7De<[f:Q8J9g:(Mfg0Gb;#I<]f=aST_/Ta<VL<=XXEI/L=IGS&>:9+PeQS
+J?YDU/O=I&.HWf=9/[a)0KS(;==J#c.US4)M/CR,)CGU?4OJS+]<ZQ=N2P32e+.
HW^7KUT0(;L&AXZT(f<b:PA(ETWBQLX89W6O_(N1g1K;9b2@:MR@YT5@1V]g]E7S
CB:</7#c(<#\Xg4L#55]g@WJ77fIZHE,U=dJ+)e141f#8-Q&C.(g2J;<-Q1P#M_D
>?OXQ]/@@U9c=P>U6E;;3@[F;YY1F8A78LaG@X3acYTP3^O#4&5X.f#0\;fIT<XR
#-=8N,4L@Vg_M9Y@1(7<L;J+[Af#e]I<]#5N@?,ABE\6R.NE5(ARDF[)[&;2Ge8N
JMRW99DGI.40I@]g6C(eAQ2F9F,D\NFBg+7d&8RQcGG.SeeCaE,_YCbWZECe/Udd
8d9a(;ge57131/+V61O/K?Q6>gLWL<Y,E(HE/;XGB(ePZObYDHD2d52[[(=fR<]d
,Q.)=/AH0IgdT]dZ56(7-6<_LeFA@;ZG,NQC4F.-^XaZ?2.0,)fZOZY3QAQf=&\8
/63IOV]MH@W-g#5U4GQg.-0fE=T37a6O/EaNH)(P77gJ,+3_T[EOcVWgEFe=&P8@
W62,]/:68Y8bD(QA?I[PbH@L=GNP>2CDWGXe[6BT]:K#K;)>Zb/&R(c_4)A(,\\g
\MFXYGE_CgAd75g6Qf?5T.dT]91Wc.W4/\-FUAKgd;<HJO)](,QZ\OY+PB-.2+ZP
4V>)>fKg#H\<,NTd.Q<G^2KD=Sg5Ka+A96R;bIM_cPK3N><TTFQM80O)3HH-LT8A
2ZNA3_V,Z&W;B\)QYU?CcM_6)W\?+#&TI:I)SQ64R1M0+W5,2^YMe1CGfgZ(EOEB
8>gH1CQ8N0Kg=:MXb,)OK9/3K>5N/=Q:/#U)PCF0S.@9)@U2Q_f,15U=.;c:06KP
^DddJTT.NGOQ6X<:-4R(eUf&))c9XE<1[g^N#MI3\b@SQ9I7MFA1;C-V8R]de:]g
?Q12IEg+,J8RcOFP.4&DW28UI\Y:P1eNR0E9ERRd2_]\d(2IHEJSF]]),2YI_?B^
a[>OA/+S/D=c\\V<We>]g(H;Ga4QWgAa?>Q[KH]2;174XTg/LQW,K)QPP-@Z@J3>
XWVDW2YcZ6HIH[d:Q\MPb;f4c1?1.D\1>U2OdQH.+?#]6F,,+dad854+BfAIe\c_
Z<F=I0.f]66fLLYG;Y;O1Pa\#PCaeJW_@a?6SW;]Ya8f&g-0e-91<^[CYHc+2U9,
M(/=.f;?DD=Ta5/]fABO5&c2>>aQARVLBLC@=&R)P;X?c\)LcP]D&A#PB2VG:;\b
O_HVCPcK?C/+(F&a.\WgSgA?c8\ZBVJ+J496.b;.fUD(deVfFf8BA?3TXV(=gbJR
60[8d,_#=^IQGF\1<O4U\)OTEOV8e6AeQX+3Q)bI]3J#^1Xd#R#/TZ\&FC5ZAN[e
,Kb;_+I,0>/gc2ffEYA^g\<V3cGG<c(R;-+GJFGb&]BH,8RSD3/0V5c4D[?aZ.Id
<]=&PF0cEc<.-.9SgU-^?QZe\)@f\GTRS5G<PPSgaS9b^E6NQ/6JFd7IVXN&WMf5
V.:47c71,^S[8JVb;ae57ACL<+8bY,LaX>1CQS<1#3BQN(.V=C\W2L)+?d/I/;P)
CXcWD^[Mc@&Y>PNO.BS^4c+b)E(00Z[c,3:R&NZ8,V2fQN2Ze/BYb]BbUDfA0-2L
.5Q1N3,[L+X8gQ5;g4)1=QH1J;AJ5?WJ1-U0)N<2M)Q/KH;>V.&fLVJ,B4H&=e02
LfEAeQdM3+9LM^K3aL3\V>W#T_FIY_.F1cO/@;8aY(\:(G5eQBE>bCB<:bMb.gQP
SOCRL]>_YP\-#AK/VQ#EO]VIbB]^7<7EF,6cH.=33.L=[8_.#BUNR_UD=K#Y[a^b
/VaaWMbCLM7:K7Z?1T1HQ>,<:1,>HZ9-G&T<RFb.?_J)4F3cg-)1>:VWg1D#bE@a
F72S:a^;XbL=JK\Tg]][J5/>e,C]2fCeORHQ^#8PD&4WPOac+];2]STE_F&/61VA
cS:HQ(1BTeMRfHIQ3\MB^NbUDQ+\A,^?eBd+3=#)AaX/MLS@H0@?cHbaE(:]X2?V
K]KU:J^g-<[d[TQTKMFJUQ)W#2.28\S^9UP\-NIX]]],X3,R.&fNAIFZ0b<Z6@R#
FW5K8?//aB,dc,K=H-+8c?BR/>d4aL-P_:6JfE#W/.-B=V;1X5MHFaLDAG.B\dad
^)J,S:7T^JVW@Q(Og>)-LV=J<YdS<^=8TR9c:?,5F5>E)aOefe.FGS7\5O_=bW6<
U3aEEf1>E>ca#<,,>7^)bKTUTK)MPBO-&).ABfOg\F)HDRO1GN;_&DIOVdR0(ZE[
L\KaEGf^W,,dD?(eV]/--UGQA,O]L89JE+SbLb>]#M@#FDG=Q[;OgDMIG^7\9-V0
[,Q1^BBc1(YIVBEDVGN+#_4D(]UB-I#d9e[\Xd4F.,QTVa-C,/431#gJ(=:YA6AU
&<_40ZK\F=YGUZ8)G@c+^I<K5&2->?IVQD;YQP.2&gRKI-g?31e\G/54)J>bMT;a
W=Q1KGZGF6CdD&e,39fT??(c7OdPA85&-L>CQU5&7-Y[,WZT(dBMWUd(=N3@_K>5
&<K&Q;(Zg>3dea;\<a_;.TFdeU#[?,)9eQV]?+YKWERQBc0NS8.d4JWE;Ib,DQ<3
_B]5>eg@X=,I#Y2HX:93=e)\Qdb1VW1CF/NUf8PX.:FW=EHAc@,\Z/e_7@:S&FK3
E2)f/BXZgbT\K=c^_L+7W:1@]IMA#]6@7/6):0T4gM)B1Me7PX^fLXBd-KVfC8H(
5U#]O>D.IcM?U13dPNe/.6RCFL22O6=Yf_HFNbB>1Bd_NQMe(G<R_0@;DRTO2WOW
Q@7b(WY?:G6J#A8bSCb=c;:HLS8(W_P>42>0C>/NF0]<75RRBOK;K8\^Sf:^]_g>
\@AO,BFV[)_=[OXV=[;BW4>2#U1LG;:_3LKd,X#cY,E7[TVB320T<.7__+E8^<BI
]OH2KT[O)J^3URE[?];cOIFM0g_c4Y@A:)O&M-<6_>.1SQ0:Y8E[f(FP\<TRg[.0
\OQEJ.OZUX3?bNdY>BC#G8#AUSQ&6N.8Z09A9M@S:^IX-fAJ38Y\d&XB>B.GE^I,
CZb(,ZaE=N5\EC+&72(V=JQSK.@./DLXa^E5@N_ZQI)ZgY2Od\_LfMA[6X)d/CZ]
18ce@@,SBGJJ2:F]5S,f=]S4cS?Rb<=\])6@C[1L;4XVV<D)ZI&EI\D5e3VD\f/?
gV92H<a-H84Z4,ONV8ecJRWZ/4B@\L,7bC],WWS7EZD;>d49Fg&9IIJ6O_R82_Yf
7=Sb6g>+OPd/JH\9K:geBfc)U;^cTZ8(:>?g\3]&aNIVW(<&:Tf&M09.G&egJe-\
SCEL,O3gU[;\Vf@8D+ZgCaCYAXO0,:7bQ(JT,WgWb&-TRQeQJT01#fg9C4g?W^:K
MP76Fe/1(cP3@M\\4FFF@Q)&5,[^QNP]6+[+M(>F]9&]AJPId)d47dL0<65B5,gN
3b2[,8(OM>F-F>+X;3^F6<V&3H]JOQ5G@PK?FW+U&L->g\A&HJL#6:,5^<R4_F/b
C.ZQ(AFO7;SSLgW,-P,D[M=39X=N5B-fP,:eGHKR[/)83dPG+B8X@b9TgTgFT;-Q
^0(+REFF-dSM,OPgZcP6PK4_+1F_SX[UT6:e5L;a:V[@&<::PN9/(_/g]gM4[M3.
2TEaA:;<O7FP:<ZTXWgE9OJ\DB9bYZ6&],>+a((O5JMgX5HI58(F6.FCW4bMDB84
:&c6:g2.fTRCcO&+W;CUF@\NT9Pcg5d/Dg4b>W7g?XU:_gO>COd^7F\^93FC:c^^
QBZ])>1/e<P0,A?>SGE<XSQD7[3-EMR[S2&KSW:641@_Q12>A<#4,P4H1c<b=E)1
-Hc<W,aZ.7H30d;SE1G85]4NCM]d:-=\@gCNJ09bZ,ARJRN_:3+NV?><3cCVOM5=
D-__G]]0d\S^bBbXY8.Ae-b(PLW,/86WH2Sd,T>WAZFF3WacPQVNUU9:_K6Q8L&&
cS(VWQXQS6KTHO9]Ma/2AW4,4C.(Z+.&B96c.EW.=R6O>.A=_C\53=VIN1B=WKd7
Sc6U;_]57PN1G>40e,c]V[,EJ<-Z[C361ATeYE@QV,W?TBb4<XIDRZ#8;>c2UP1.
,N(<F,)=)e+eBOKdBW/&B4(U8c5-c9ZX5<;KI(gCRW^Z1?K9-Q[/RB)_NR6BO;/F
@1IaPD/5?Y>FBRFJb9Y^WCbA.]FN:)]<50a.TO+G\&=B-YQRH8Ie5DX08+SU2FS/
BFIWG<+UV&0&^U3E<=[\GJENHG2FX<9;SKX,PaQA\(T5fS2E?07IR<R=RU3F74[e
P,V:ZSf:AFNFU;;cX<./0GeHX0@3>[W3f_[ASbT[S<AJJ<aC;W3aHa,-Q:gC/,U:
&Md2TMeRfPRRI:P;N6VTgc<;#3L7EGC0FY@cDG^[D<?c_dB9aG@WG,-1;_RJYRLI
?@-]3LY1O&X7>QZ^E00\6[_[=E?,MfSW0FE?:CPbP;Ce&(dNVY.B]Wf:@[H/f<4T
=F=QWY(9)4d.FXR>J:3_aaXPM8WWJ,+X_\=-E/WNOMIMEAO5?D06&1Ned@b6Bc]K
J)DRcC0P^K&9./YBge\>+?Q,SQ+.Xe\X3DUV]-..Y-]6?;VZXbF=+C)TFJA;>#d-
@)C1?VAbU/g@)[=)XP<]RfI@C:f;R5:PUEKU<c>KWUage#IH4#BEMQT20I>fa,EI
\62;>5^=)&Y<4DF5=Ie):)21H9\JP2QgYaE-[).C;KPa1?bN,M^NO\/(J^CE_GHJ
]2gU:V,PLN5Z;eMMNa#/4#X<93g<]P#cLC/_4OWc+E2YC8/gULZ;N:d+=XX4=a19
4S8)I&.e(gAD[/33]I,1K)KSA]V.D+Gg_aR+4E#_6cO]3Ub;g[Y:SR5(@#;V##Af
7PK^gAMQMeS^=<,;JgI#>c6HTBF3Y5H-B<X@CJ)WOC1aXVae=E>HAPRO:2eWF).J
X6&1.0@<eYa(17-7Q(D1/L1I2UD]KF00=I-WOR,FB([BbTGZ&RF6E.IC.G9>3<-=
FQ9E6.KIa;[,+0]MV&RZ^>5aQLH.MN^[gJ\#/+T+E76f?A#Q.^dN>E/+12V:<IEI
_.M(P2U7=,^Y.5E,Qd_VC&Z.e8[GY4<@INRHXAG)@bJ?9;8bc..c+[^(GXe[?J>9
b<DE>IYYBP+KUIL-]ZdaVF,@3LKgCP30d&f>@?.M9TNREOW3(C5PH2;.P5c5?+cF
BSJP-2ZRF2LTeZO_b=I<?@8#,BC.I;&+#(X)X3&NQ<9QAHI1IKQ72P@DVL;M,\4Y
aXa(SZf4^cVG,dZDN<5TbRMGH7T/GPH1.2T?O9PAA[A4b/)7;Y;[HfP??2;5NeS8
.cA]KQW,-+&;._M+/fJ)D+HEP:0]&8HbH\-K@VHZHgXIAOdQ5&&N:>JI?+V/FGTE
OSa2?MBLQSCT;/-(X<U36MQ0<,FNBWZgWa#HgL:O=a9D.aM1gSOJ,A3^:_^P+b,4
FT>@P1AGXDX52?R]@W>I40JVH@]/,\K;?3->\=Y3#JOK5@T7OCdYV5b6d,Z+-4Y.
S.C0G@0A:RMW?;&E2(8@J1>gRa,+[g2WO/;,](:X4[;#P+a@6eST&A5g8:)0.O?b
_acJZ;9Ma(Bd[]?9)bMNXef_MN@FQWE:^4R0)CSNH##HHURG[SGJaE4-/XMU;Z#C
;JYI<0&>J6F,+YHP=8VAS,>g62QJY0G73[<NZKVgP0O1dI6S1\.)C&F=/B@A]>PP
76b;8D>ZR(#Z9&aXZEQ8[2fY;3@.8e7U:L/RIV(e>3f+d.TP^:L7XGP4^IggY;Ga
6?eZg2)0RX_E+3/AgPWBH;B1PQ@]DSQRZ?S+7I#>04bI<Rc^QW_S:9E77,5Q7LP0
,)2,c#/d(>c#(e5@#DgKU+#fXf;Vd<D(O,5,<U1<CEOJ;Y#DPNF=8\dJ5,^_@(Y[
]gc3ZUEd]8,O]:&>WYFXH<F@ab?c9)@,0V13ZOIUDK:9Wa)UP40/E\[JEFC>>D6M
eTB8581FgAW?f38W\BMXP?@+f9(aLL0S?@Ceg/[\WG;@K@E_)UUA,IZ>YR[1AeN3
S?9P-QIb0UQNC?@>aJ3Ve:RPa^9^)?N_T)^/_7B>.HQ.&@c_KJ1d51.&S8f+^+Xg
.RXeY_-_gW_4S&fUG519JFODD-]LJ9\)QRKdP\9NPL1&TI0<@?M[B&a:_372&6K0
cA1LP)1ZC7;Z/aFZU9U/(P</(:SR<+>0cY44T1Oc0,e+UIB^/[J5GBK?/T[P\_<?
-JQ#^KNL9_ePFV>4E\._MgIPg[BWc5(NRR/,/9SUK:VD^b/83EI,@-1(H;;:;[+Q
#820^:YR9\E87+eD_R8Q,TfF.Jgd6L@[CA4XBS>cXC^eHJ>8d-(#=&6EA]dS,_O&
F>_664,g)@]E?AIC>^=eb;P[H_;#J9>FU5W5fPJ&)cE6Q9#HC;3H(E9;fE.DAJc2
B8R3XH>86?C^?W]RZ,:?D,d#U;Nad3#:^URNVfMAE-Z(KO(HG&O:gJDc-e)K.P+9
EJSZ_U.F;1M62CAL=TbA[G4F1X)IbZT7)K:9CcX6EDY2U\:EW,.9#R:PNUBN6&E[
U[UD/g3_GgG1.03]ScfYP6C<M4;@;RIM5TAKJJXP))c_<LP19-8FP_QDb4,,cO#6
A-7AUVY>][E/.?C7)VB]2aZ[GK:VdH.Z,R]faRDUaD(fH:M\R6(TOQb9)6#[M[3X
N,=.DL3@35M:N=XA9FTQeMaU&\K/_>bNJ6b8^G@IFaW)KEY5IeR-gI=DL4/3ZL/Y
OZ0K>Y5_=RC)UUbZR4cMQ)(2XTEUUS/2_O+:N.Uf7=#]f)5J=A(-5#OLc7cK)Q,D
:AR#?/2,L;@WXBO>]MJI6S,:S86DOcMNd6MbaGc#Bc/H^T9]5]H-g/BdL^Cgg=/]
-I1;PI0<</:S+FRYD-7)5_GV):;J:]?^5XU\/_T-^#Q>AGH/;:Z?c4-P;A:_D?@Q
/]^dgEO[P\K\&9d^SG,g?>,GG+9bbd0?W<DMT?H3624P_Nd/D,M)eA:e6#ETc61D
R7HFW:c)9Te<[H,=7LSKR8Cdf&1<H]KH./RdL8[/=[ZSOJT/F[ggB8/.Z[XJfLFY
XE/fWBRGO;NY\P1VHR.4DO:,[\3H?C<d((.g5?Cd[E;_.e08?,8-IcJZFdYA?aLG
G&XfY=NNEMQ-_NWDSZb@OHdQ,>d9MHD+^C_.C@c<@C>NL7Zf^XgIL:TZ_?Ae#M3;
GN]:II:A:-MY[Ac[f;>aH#NaY+6@](D&Rc]c]QXJYg3>22[eUFQP-.a?c[BcUIO8
XVCdP2(98A:VJDN<-,AOQT?&3cAE:b7;(,#0a@.(V<AI(gHA;RM\D0.MP2fFHcZ,
S-N1PO0f;6gHP;Ec+?:Z\&f/>EQI74?@1XaXUWJdBe;c3Hgf5BWZddf?;RTEbY[;
C/ECU)c;aB+&]8BFC6N4U&Mc<5[:[)V;:8,X.7g8Hfd8,GQKaHPK&F)KR^,ZI@P9
K\HgDW1]SKF@B^M(_+Ga[DE1>=dE?gb4S<KRGO+]5Z+C\7_:U#gQ#4gg9T103Q/A
8&JXPR-LLS1L5&fEN[OKR/40RbX/ZY+W]e([+9D?&.&TF5:S43I]dM1P4W#+A_e/
#OaAGV>_<\4G43M[]Q.TIg;^]c(,)1eJHY&05MD[&MLIgFAf[MNc+=:C8I.MP8IU
DQd>#V@cZ)EH^WF#&XDJW5WcYE=#<TKX2#&ad-(W2<>dCXLC\f]f>ZCe5QR#M:_Z
.Qe[[A;.LLN#b)VGII?NMfB>:5La>P(]]b5IgV[1;BV,@40\YSIN7&ce/>RUJMB;
=M:K_PSK0?A2KQ@JU8Zg=LY@;C)9F7ggf:OSg<>f@C4P;U?8OP6R#a;LI:99U+^I
6fM=)3<;-C1f<S=]#4+/9T.EBA[aQH5W@gg[^74>&2R46K3Q60S&H,e^3^.OKA\g
K+CJ[NbNgFLDX18#.#O[_QY(GE7^:PDSQLTN:OHcYPYAb(GR<6d=7,G;]R)[BMA<
L9RB1cO4?OA)Ng/XSO=MK^Ug6ZNW<bf:8a1dP1Z1XeQLKBb<47+L2[IMKSaGN?L<
I2cAD6:CfGaPZdSRL4A>+ABZMY15NdEb-N?ZG3@VUX:JFL1fD71NQB\OF:Z1H)00
3-IYC#AM53R:P7LbNEc>/d92?9.dHeLX\UT.DKU+C3CM?28^CM+Y>[UCc@HS&<[^
c6=f15BeH^dg+4W\J^M(3NLD;Pb015-[MP-IA[2W+G4c[PE5QI1H/L6g_T#.gER7
H(A9HMd3(d;J1LMb:bR5EWZg0:=#R<g4<+=&EJ528YZM,TEbOI0]#]R5O);8#QYS
&MRF;5Y)+MT7&A_I-6DIGW-dLaTJ]W;&(BV<(Pc8,d3=<HcW#LEaTSaRZObb3?W=
OQEPdIF\_fbbY&Q3V\fQ@Pb7/.FAYOO7Z\RHLCR_U\(cLf3+BKG(B,]72X)LLX7_
=\X:VGV1c-A-5.)NBC6#5(Z[SDYHE<?_\Gcg:JHND9(Db)GS/;OMQ^H.cJ7+<HaB
<>KUP:B.SK=,QPPW;DfF<#KTCT]<+@X1@=#d2+@.4Z9ID;MHXB_INH^[VC6Z]0D+
I.2T_,SI0g05H#9+E;EB;CAZX7]f9?[f9BD?3\=+<?G3aIQc=&X(WC-;77ER07CM
S#4/cP10^B)>HT=T)6,+QQ+2=<IJ:V+9a3Sdf5efA3\c/Y<XT=1[GF[aD;19&C7R
P\f80cSY.ZO;a3a_e8B_c7c^_U=I4Q9gAJGD6EV74gg(C4S-NZKA[WE.:/3W;JXI
U#<;7/e_53GV0H23[]VG7VKBa,3dIgBLb5Ra[0P:f6B[F\X>gH)GCB^SDeI-]dM[
FQCf5V-TM@PQ<bTF&b_7-GO(@/fOOO/X+L-&\B\T,O/<&IAd<NX9]gcCc)BR5VEP
3b@H)4;1Gc\_(Tc2XU\31-I?3_WFX8e.BIc;ddcZGeQSRN#c52/8GINEQ3dBWcAZ
CWfY5Y3[VQRA)J^L6B<WE.#CdWcR(30dYCL)K]8YCJHP&;b;94N^VKHLeLf@S&OO
#91H)eL;EWfAE4+4/9=gcT0#E3^:2^b.&&8;2O(<:8YABX7YJQ^6A60Ie,d9g9=c
PD4)Fc.TR?F6GM[9<^APe.\PJ?QY5#64H3_8e&_bc[W,:&Wc@,fF^f?YH@Q17^OK
BF3#eW)#RA<M<#H<J6_@\#+X&AVg&-JYNXR>=]X(a)[SE]bS0b+3aVU^Sga1G00f
M:S4GN1EP&bcMS2[0\.&Qb8aKKD):H1N/QZ:H[aV.=H^L&CdG[\fTNBS?G81<P5I
.&.f#eW2T]@efF3?R.HaPZV^>(G1JTB+@ID[.IU\)aFc_I4X&([[NL/]Wg/UBM6B
^O@732;g>-0^YMedC-8;_#SHR\^g;bRDA:0^Ga#5\]aDG2bB2PdC_CgFQ5((De/^
;7-WaWV])L-ZP#3f6<S7g3T]QK2-0_0)XcbR-I3NUB_T<W03G<5A9F7VM,8-dY@;
1T024Df/5<8/166SgN.U&f1RD)AS8\:U-6c)4;?2=1af9aeB3/5A@;g:aXW>GdWC
^2=&(e#BTT1?64A)g4FWW_RcS9eW)3^J8L51I5LI6a0S,)(V9:a1N8fO<51M7.b8
GNSN;O3>9MNPZE-?RbQ?6MH#E]ML<5cfKEMVfTFC79C+.2:?B^R_B12#7^B7a1Zc
H;\=.0BfIC&T:@ebL-QRZ.6;YP_Ka;A,fU\8<Ec3@SJJK9K5E6e]X)\\fb42C@5.
0a/_LZ,0-B^0=bJ,>0ZGF:d#FT^:JVT,84:?(>B2^#FPc(NZ]F9N)c:?8+/WZW07
05LPS2/:>I:,-Q@]PZ,@dX&8eL>7UEDVa&DSJ[Y^-SE:GM0?5eZHK[bVKGcJ#]30
3TA;&434<e/Y93&1g/GS^?7&_MO+D@?O7KCJCKF(QJJ)(.)NSNd?@XH0SQ3A(0NL
8KRY+>YHUTT2[\c19PH_M^X8F<dHX93?=ZS7_g0a?FNA0=E[2>ECCT[_)Tg1dbd1
]LSNdAO?^(DF-e=BG)-ZZJ2RO(19#b2Q\+)&eA+@V3SFa?3Mc-)I##/3UEcYf=BZ
N5@7JBMc0]<=4R3ZV2<_^^B])CcS)C-:,Id058U^CYXPdOX6=JCPE,,X]:Ne9D[S
<2e/Z)Hb+LB9+/AOS2_HD-fA+)HC=@cXMdS4\MKXNcOfdOWJ49J-D/e<<_8#9@AQ
eK)J.Z(\HAX^&T2LB22V1&ODFD1UO?b]a1&7\7J?U6#Y<b8?0f=,28_W8I?YVY8c
G+9IJLFEe,MX]LAH=S3/Qa)LE)5NKXK5YP/R6]1L0)[+,)W8AS+BFF135OW\CLL>
ffdg>EIYP\69W,YB67QJ;F5c>e<c7\Y5ML)5D=-eA(+7-/]Nfb_H<[HUDT;PU1G+
J8bZIJd/d&U)DX+9fe>OZ;TR/#P0>A(2G,_B+#F&I(0-^FU(VNB.YP)D<5\(01&#
M_BU[M:)S0W0.)QU)XP3d,&Qd;QO/BWec.H<O_^D\f?H6).CgU;S1>W&=JSHY?GW
##R[SB<.9Q4@CXUQD>QS<\POAg+@:gZPd:YE:?0YS?A/B,2L3H#Aa4CHB:BBJXYR
=>\Zf6Z.<0UEd4O@FWGXdA(35egOWE4Z+JObU=LEF@AW\]+c.0-AQX5Xa=^Z/5\Z
#;IEX3JQ<D?,c8WGJ&/AA-2AaOJ7G8edRRdSG)Y#2#0]03MB8EY]B^S+5#B\ZG.4
e+;HG;EQbUUgJe]WL9<96LSY]T+\CY[.7UCW_A^@:7JV+I5#9J@B3C/S&d\YGBM]
?\c,a=abU5XB?-0K>:V+RPaX<312S,G1_\P:I?T@X67OHW3PJ^,&V4^952^e#1=S
=UFQGAYUWe@7#KO(SNX\4G@Ed[7_8ZGdTI^#^L4f6IAE9c^-,[VGXXFM=P1C)a/G
=XP.IZW3c&2aT05IZ_\bW43QeN^4+d&##7]QAf_7EQ^Q+KV[C8GX4K)CBSS>(7<U
[@:9f,CB37^9_3L/(F4O_FcV9E1-K<I@\(YW&=I00.+A8e_^]HQ(E40c.U?ZI#9<
@#SF5Xd9V2O?00bJKVc_N3TP,@Y:TS.TN3V&);d0F^U7T?\Af&TgQ:=FZ>>90DE@
DBId1Wd@1^BTK0XLP9NcB[\)B#M=dg&Y6g;V@X>)NH,.>3+>E?@9/9.4N@HLJDO.
2#T]QG9AUQ&APKOTVf1>c_]E6DZ.49M7[<MV_HP:=D8XT8)3CNd-X>IHP_3gZ@\4
]HNa(PBBUJIfHN2UM,:.?5)J)ZD/;Sf;:)EaN#PYHPGC=F]S@HNaG8f0#Y<K;3YK
16S<CFM,_SUb8d4^[.Q6C\3<_F&Y1R,CHX.(4?57-&4:RQWfFbNAZZWLIUE/)W0e
;4.\0U4/F0=@95aa]6TZN<1US\0TNZX(PMXB^Y(E=:=2EJ0:fE\IW\,0SE5g6YUM
OW4c+Zd7)Xc@ZaD?b#@._Y9(>[@f5,FF2J&E?cE+c4AHR4MgVcaKeN39+.H#&YF^
?PNR;B/aM-F->.W0c>C,N8[J.Jd)NZMa=aIYQX@c&QVY_(PCN/55DOG46#g_SWK\
Tag4,B)_/2d\G@:]D@aAZ[<RWPUaEPZJ=CA.](Zd5g?dfL7B?.:I93W9/R;8QU44
:\cPSB)LD4WL9d8DFFI1&?75-7VM,AB?;@3BJgH9\>WYJEXICLF\e3JL?K08D:E/
XR\b7Ng/L&N#9:I4TdgDY;-QF3WR)Lb,5bA,9P:N0cKINT[N/X.<SK-6FQa,A7+?
bN.@Z-K8LBA[\<+:W)]^[S[f(dbLdN3YC.\HB]3>F49:.X5PL,,HZT#9DNUPEC=[
5M;S=/BVU.e4^^\WX0IdR5d599>EO:5)UDVAIcL)F8=Z4JW&NZ_.F5[KDeM@a1V\
Uc(L,Q)2GQOHYZK@a(Y][#A&STW3W<M_+,:=/a-:d=,f6FV=U:YC-=EJEAMR^:Z\
ML/H9:@&1;002M@W=L].7aDQBKW7ceFR/;=Ta_2Y<5V4TO-Y&P7,a9Y+9H/aO309
FHH&9^Z]KK5c]DW9@,KVB-AJ]-TcHX>SFONIQ-?94_E&KX#HbQ(<IM>b(eOBc]+(
LC>NC]W@-LONN?C&^7CfR8LY@aGMDFPHMbH.f7ZH+bJ&LIF8HHO]Ed7@5-2W)938
^G9-QR30Pe6g4b4_/EVCOI0DcJL?ObKK)+Ne/7QS.:F,3C()FG,G@,f8&EHG(6gB
WUE@#E#S7H_UeWX9DJ)S1LPCR#^8JPQdBaC]M50->5UOIXaKB@FED#=5T>TH@_1;
7Za95DX1F4f:4#4AT3J.388&YbA_>Y,T/^A79ebdb5d#D+OI&bRcA]NDY<U\?K(I
=K-fH:E9?M/@KDXSL-F_1^e7M:8:3bZf>(3F+d#a&:@c7GSP92_;d+5\W7./)THQ
2154H-Y,TXcDI:U,)+ZIO<Gf@]V,fQ(.0X=f-1.aJC&0,Z:]:faUM]\1A5VA(GT^
?UKfA1:K9G^85/_B8X?BGB@Q2+]-YFV@F-LL.b:DP#QcSP#CP-@c<GH:fXTI-K?R
MNR61D(dSO<TL15\WfV2^PLZ[b#MgegFF\L&G;BE6RV<).NEE;.#g<=XMU7&O_V]
MZX28bZ\D1KLVf+H1JO8:^,.7/Y3@^dNX6V7L/4FO5TEY4BMQbCEZE,>E5)(+\,5
@SW,O/UQKc+3,GX[2>A#)Z.,dN,^0a6QGg@_VI852]CTUKF9b(K_4_7A5g)SLDUA
]\0Ia;8T[:Se;X28S6;U/^ZL#:IN2DP[H#=3C<QC&B)=e-07]=#IR(1g0gIEB[F6
gL]NRA8MD99]L.MSGfL@/^S00MS_W@_?-G[8;dLV^=H>9@6fV=KH5W]X)X?@7V2V
#N=F#,PNM0UL5RUa#VMJ5UY[TD<X#UMC]@6=^#dC+L5/#09b+Y+EY]a,JRCG+(37
WJ1<_:9HU[\_gB/7(?18\^Aa=9XMg5\H\BIKVTM;HZcgTe+gW\LCRGKfH/W-,4O)
I#AgdJS2eB>F\EJe:3Z8Bf.;8ATWeZ;YE5+HZ_(3++//0ZggDWXb(77ART&<^A&P
7-;bFQY9KSWXVG),0<g#.[9,]1-DQeOX3,]L(_,F810Na2/54U]Z(^g/-CF[W(U<
]H+ARdB1MDX.\NU_J>1D\,aR7@M+c0K7LZ-+gC<9H#K4Q#SK.T+P1.59SLW_R3,W
eeb(QY-2#>UTH,cX#;@]0S6D)>\c.CU+IIXEYAE/JM19,D_WQ;,<2g#MfL8Q>Z,H
WePT[-3b+JdgL709+fP2(VY6M.fbga9-G>:OZd0-DVBg^\8>MEDG)Jf3LR/T[:<K
YK=UUeQT]@)(^OX_e1gS/B)Cgbg?V+28^^&Zf]20UF13bcM1B2;<CeAb.V_QAfIc
MGPRaIa:6dR:A-V4(?dN3E#)83PO-2X&]252>-V6D:aEH<6Te8+gUNfA>/)Z;WM=
OV4R2#;HG349Oe=Z,DfE</8c^\a(G:@Z>\([_:N9b2Z&-?]?HNb?Zga?;_>F;:-\
:S09e3]:;d/Cfe&6H]f<\STQag(BH.S8)/O<(ZVQ\?X02>Q,07NB+UI-<e+N(dUA
#I,J41Y>EH-&PM)B4K0I68IIH1FAIF9bc:O@B7:bW#6Xa7(O1.AJ3M.I(VJ(RHd[
.3^<+:(3g&eG.PQ.DRPX0Pb3.31<&d)(=Y@eR>&:0eGa\#WH5K3LV]dP@[cA^2NK
9ccOc_2E<C\e;Z#/Ee-PW.SJF8/#N&T2@JM;bA&[Ggeg:-;eV<,1_,(:\cI8KO:&
H:G.dI.M7NNA6/5&)KL41cJMR_L]3+IW,5IP9f_>S4WQGN(90,,DEg64G)BQ7/]E
L?LOTR4)J.G<)@[I[VBDFBW=N]9:eH:]6_F)TD4-VS)51;]U2>TO:;(O_JS0>Y2Z
6W#RKZ+)f[1YGX[XVKdJVEFe0KU@QRfOV(fAM_ZUQeeW>C4b+,]OVNS(LIaKOU/g
7W@NO37.g>Ud.?ZWfLLJ-9BUd=-OB]#=IF5X/e\\[B@F#=VU>d/aXC_:b,;,9[G#
5+0UbcP#b9d8EI(HFJGb?YdSJSD[6SPEISN<Y>\^gFL,,><b.-0ZIY1_5YWAgD>0
T>-VNUR)K],,HG@ae_#Z7HN7\LH3U@0^Y,De0V]0Q6]<P,3[4-H[7,.Z_.D^e+S)
X?09McH^RIR;BM.WbcY@5>]]g:->_7F<4C@IUJ??VfQP7J/)eG32b,<[<\53(^MY
P&VBX]_2O>VWSbFP63#H.GVJ31.[,N^PDg0KTH:gTD,=c>Ng&#gUVNdc1UDPZ[>J
dRa40L(R>PY;eG/L5GA1;OH727#,7&P,f&VNLEE/@\dWX0gW4FCB3ReOAfO3[>:D
H.4:Z/L>D&AbT.<N&QVCe)FX:b5YX@]Le>c@SFX_d2Z=VNS-f007S9=RR-BM[A_d
@LBX&FG;YXQ>e9].Z@L4][L&(+ZJP[aCCXX3[1<1[)U=1d7E4LKC(()N4Z2&VZ0,
#XNbIN^S]E4_RM=._T54BGbR1GHN>a3;2X67CR_d;CGTEI4g6cD+I6/S>#WM:[UG
>PS=#&CL9bb-LI+GY3F&c_R?dMe13S:L4Q4-2@QH#6)B)Xa]?0]XZdA5YJ59+D#1
aX>].&5NU<HN5.fRX.HZH.<71\[LR)E&HC22JXOPN42bd2c4?G.;EG:145P/KQ^,
78<2CQG?7f6U./UL8FB+<F2RC/H=2P\[62:9B58d0Qg=11=X]MKfg.2TWCc28>]C
1NL9+J6UEMU7#NA0B?VOVC#,2YYI>3]MeC<1(a_8d#2<IV,E,\DQQ#2(#(?2A&YO
O3C63XKR1+N.-W(0BeQPUQ_<J8M;.N+A9$
`endprotected
