// TA demo pattern

//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Siamese Neural Network
//   Author     		: Jia-Yu Lee (maggie8905121@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      70.0
`define SEED_NUMBER     28825252
`define PATTERN_NUMBER 100

module PATTERN(
    //Output Port
    clk,
    rst_n,
    cg_en,
    in_valid,
    Img,
    Kernel,
	Weight,
    Opt,
    //Input Port
    out_valid,
    out
    );


`protected
41>R/4[:Oa:4dgS7)4&CHHL@,9TKXP=3EO61a<YcMPUV;ECg)bS8()>U(VIVO0(8
e(M?H7UAa[(Z=M+S(fVBQWAK_D?a&UWKNQA?XAM(9[,ac+6HHXH6R<HQLPgH8=24
C?B]^beYb?bV>62FOcZA.ag4-OH7M_ef2_ZX;GGRa<X36WQbT^-CgOe--NZ^17-C
[-/W4^-d..+O=L@4E?c^d-5K4(I=@^/<TR74=MO(=@H(JX2dXZEJVCT5AG00=H#O
GKYR0\fe:dG./[8]4JK)<SGMeT<d6?B3=#PEaOC,^9Y?OO^<f5@06>T5K$
`endprotected
output          clk, rst_n, in_valid;
output  reg         cg_en;
output  [31:0]  Img;
output  [31:0]  Kernel;
output  [31:0]  Weight;
output  [ 1:0]  Opt;
input           out_valid;
input   [31:0]  out;


`protected
@[\9Ca?aBEQG/<[7S6BUNOe;<87QN9VfKfCF8SKG,dIcW<b_g2WR.)J#-^X;KK?7
53W7^\@GEf0N9-&g^Y9^aD1E(/X^>)W:LD(9^06F+_;2KY7J1>KS]-DS0G+166=6
>bIEb8.U-:@+M3b;/Q52.]//IPF8#Z@LXU+[fc@J4SIcK6,Gg1]Y)b?Z>)=V@_:f
KegP\RPAS8])LW=P;1B[B7D_1Qe>[&R1KPG&;gdDWdUK,LHGWeM=J[A<3ZX>0YXW
CRegOXgOZKNfEdYWf,E14f58BC46a48.3e?A=W>ffHWbJ>/fYQGH)H7.6T-I)]=V
S3YC4\-E)R9K.GcXReW60;e6^d(3fNJ+XGH[Rf=Wdd)7P1aYMWPaD[_>g>&LbLRU
+4P@W3)P6RRCf=_Q?f;6+D[.ET(X4Sb]0IZQ=fG=14KQA:0\6CBUeC0&8)U4BY9Y
g?+SIbZ]2=T)3Ib@K-#4NGBbe4K/e6[H6>c>B#NZF.b4G/\:_4AW#_P@@1,^fTF:
9f(RXHA2TQ]<1)EObS(=>&8F[ET?O(I5:AJ<_JK3UVNZ\4>8<]\gdS5_=1NZ:3WB
+;_KdUQ;.Ic+#_SRMLLE^e^F=F\e4P-]eVZ9OY]b(H>:^<].P-3PV<?Wf6K_gSO0
d?OG2[9P=+)SN.LRSZ6)JTUaXK;aEZT3Me&F1-ML<M1#-d?Z;:<5_NCF=?.&QE/?
\(H(XC^+\X9>F3_G/PPRO#>@E^b,cf^5O5fFM9a./@IYY2AaV6?4I]=^g,DT[(7<
[2K]EfO^#</P<V#.4YKcQ@:.=?MXA^Jd=bVeH-f\Q3NJScSDZ4K/4T.TIN\4P/##
6[gNRW_aB2L<-eD8&Tc6981Nd=_NZY^<fLf#F@4:,:ZA>WceK>^@EV^e&CO&:)F2
)5T8EQE=4&#HM[(XdOfd3_H([YJg&dFcF6VA?V^_Yb#&O?[OPVZ3e(0:A(HCO3T5
28EW):@9]gT-gE\fR=ad@WTK_;9\NW_.,7H=(d..U^J9?WgV5E]HPIJS[B(9SR5^
eTHdJX/V9a6?]TWO7Ua5&&3^Zgg</[?0<D7/?afTBI^QgJ+Be>EcD2/g=6+U](()
8=)LMC<A2C]4QW98cO-,EAO60A.V[?dLRd5.,G39XVaW;@/+We1L,X#B)a5a^Y.D
@4QbEe1E4&O/,46M406Y@(:WCKaYeM1G#MJOK?\PSHKP8B,[1#[V[CFIN)cD3R(a
FY4A(P@3AG=aW7&@B7X<#<2K4JD<T3aWf2]^@,.Y3e[dC\g6E0:YdaOgU+b97[05
3I2gXR:V>TUJIO36>:.S?4XG3.@34UIg,C<FK2@;;dDRC16,-HSB[R4A-HOgJ0dC
JdC;/Je)GaEBVOY_^3Y/G#:>K:3S#K(Y[.V^N1G^LdOITc8E[Cg6aJ8F>c,QK>4U
.,5UY8)BM\9TC>LZZIP_f;P&=\&/3V;ORa-I>7;cS;Xf:O1]N=:X.XC247PaOBT8
8A&)UIU^0T4S>;FP/aZJ7&1U,@+;g+_+>7ILFB++1]8bXOO><FU\0a)Ia4UE_5dE
T+-B&K3b/9K@QX>KF,>-V+gW]@G+(W@#f\IYBA#RPf9C0RAR[IOY2/Db0ASgKGI1
/@R-dF=TAO_&N&]6_CP\Pc9,bX]8]F]SI41JgNQ_216/\M9bGZM+[ROYEF]QQX^6
DB9cQ@?>O4SZb1D4\(U&3aF#G:cLA^d93))KRg-_MIS&WK90F@_&7\]Z&JM8ec1:
3VCE25&^7ZI=/;_=++cX30@5:^=[:BBZ>N8^=FYXN1:7=]BcG\;^_2=?(ELaZI8V
a+^QUBeC,0V^U716.F3c>[X^PMb4]3\]&GU1/JG]O@IZ/-C9G:;;1fJ:K4a^02OH
62M[c3QR^?A:T\RG[2aRLbe4@CQ-@)NJ_eSR-EFG]2SgM,<5I8GZ4OBQQ1?A-(B0
De[>:XG<N\#IB(GY?c.S#HW=(RTf0;g6D(<EU<&2GSL/=>V\b^dE)&>W6EHZ:>eM
J,.@KHBGJ6DR_M-WcedN^4CDSUJ)Nb+f6:9-7:f/bG4YQD>d4=,3N+GN>LRG8WB4
ZPJQI49YJe[[^QHf5gP]:/00<PGYZJ22)WbcFC=a/CW,CXE6D9>1C)G9Zc=,,_,a
d3IK-CVV0T@:NOT^5^8NCQ\U6K&8fL).KfRaQ9dA9^-UU&^0I=c:XXJa(U:6<=Md
/Z[M=RUX;1C,gQ+gN=1bBMZFbNAN5MDM6N5d/5W?3>e-+b4//LcZI0<]SS]A]&Yd
<B)gDUEfc0/;;5=?]DA1feQ7A0<S(]X<N0@I[F]60Wd7X:X<]Cba;VSe;U<</G\6
cBVAII4Kc.=_687UUUfL;EYJ7S\ZT5N_I8^QE24=WEeLG)U=GG2Qe)E+5cF3K_N_
(-YCAL(IYdD5c8O_:g;CL&c#6.DbG9Hg;1E8:]=XW8?B+&.J/FUB[W:&.TL<-4YN
A?86+IK1+ON,;V\bZ#Va@VLX5DgOA2R941E)B5V[>6]=;F1B+^91BF5:Nff]U9IC
M-d41D[7FVKG]4CXN]:Y?]^cf))(H5CVLF?3&R]D@YGVR5N5HVBU#-VXd>.b(ac+
aT&bJN2KX4-BfPa\BS.)gA^&cG:0PT59fUEOC_LYN9;ZU/@6>UPL;WJ;a90&H+&2
)<-L@B&WR6)F+>Ag<M[7fZde9a7R<3;d91<_2UW=UQa^=M(J.bMQQ5:\>Jb+B#Y0
EfEFJ&9K\4F)fKP+c0Tb4-Rf9OG2Db[UGDJgIZBeUPe,1JD&+RUG:4^/-E5@ZC_X
c@b=W-Q?W\DO9#1f7YIZY-f/AA_LU]OR9FMF:LBfLUcZ#9:Y9IF_407NfM4O^90=
S\JTaR)3G\1TSR^UOR7Aa&PWbGeaBSH2/\E1(N[P^aLC/1g)NZI62)ON):A\Yg_=
9^-X-MLH/RS^XZ<RB-LTN?V:7)_L5<V1[ac[_bU2Hb#R+JXM?M&BOQ^?.A]O@VQ\
G_#D@F?UW68=ZLac<N_NU[;f]<R1KfZG#E3#f08e;[X>CbT9I99HMRa;MZCW#+g=
HB&:P7)cM(fE/cKOR0GX(^)IL&HBe+Gf^MKQ^+0WX3([K.2:#cG+SH8J(afBGc;b
aA?IPNE67J0T,@^2300:]3:8W_Pg:ST/A<ADeSECd[c[<eG0R=8W<CL6S;)<CJgU
]@\P7f?_RRTcGA+f0()Ef-,S@<g_4E1IaZ(4MIb1_IS^#Dd))O&c<X)J+N7>[I?Z
Dg=7\[M8=1#ZM3Y1:]:LWG8IZYCX0\48XKNR+4^a=VWa(&4VC9WgY6ZeQY]P2N>_
0/V<\1[b&TU=^J@e5T.0&Zf0TLN7?.Cf\)5@b>cITP0KgXf5g(C;@MM.^OM]I]6N
5E8ZN0G]TG.3gJ4Q6N5eR];M>Z5T,T[BO8J9_YV1VW+YP]^RD;[Q&[G4&f6a(KOL
IM;dI3I8##9019QAE,T-;64:C4U.M],,6b7X^TVIG)47O^gTSXH_L^7KI55Pd6TB
-PHg@@g&Q,1YbUVaTG;M<B,C8cab1Y<^e7\K0(:4bHC^N):5BQR2b6fUZQW+eF25
2.Wb.+0SFU(ZZF#9ANEDe]LP7RB8H[KIS+KBLf15;.X)7P.]81D:Rf\#fMT&19;E
-9aWBH=@IbNL2;,3)]&&=7+<))MAb.]9LR<@dad58>HgR:6>6RDZ,7;7.8NVK&IW
7b:3ZZ<=J#K6cUM&_X9Ec\F\.9UKZ^]6#C#:Cc4LDX,8+05?a6QQfI]D2.?U-HB0
L\#0<<cYOQE?ffg;2b)WgQedOFU9Vc#C]2CQ.VYY?a8VOL-RSB@F1R.8Y3@<D,B6
?]AJdL(a=1GS5H-^gUB2ZHSB<d4(7LO>2;K/O>S3<HRZR?Hgg:I.I+SFB\RQHRT/
DI2/<0:XV94P#dd0g,_Ne[Q&46_9YYM1H.-W76&@LQ3]:NSR,1XHCfH36,@<V1@_
I@M3,9KL<eDfCeGS\7:PX@C<(1T1)NXL54H4gT^II4^_He^PXe;G]#UPHV?Wa[]S
<(b,QR:JL.9W1-D.=7/K[TV(^C(94)\&&WEA+5^CA988.C5N^>WYdV_b6\\_8VM@
DA7B-K3,5QI1K4:c&UMe)dL,[V4&e2F,NG=Eg?,KJP.TB6/La4U,gAN-,Y^K42?)
,G-_ORGa(9<ZK..a6@36:+e<?d.EUTd:V4.0E[OG-I=:\KVbcG0H.:,^[GBS?B>_
-\\C5f\>R(eBAaH)0U?gOEeZNWS?XKYMN,^QdY[WaSGWfVST@7LKX6R#E[^]X_L#
E<15L?WW3^+S#7.7ZEdEQa.]PN+8+4@a0)9EJ/?P&<:gPC+-_b^68g@U]@J?=(Q1
Vd/7:?\/V-Q4GAaC>4>NNZ@<(UPX;b2[QL3A/N&J[J9f.S]84.P1-E,H[.Bc#\AH
G\XgR_?7#(\LT0]O:5_+0Q;5,cIP#(A8#cF;9N9]H8ee7-R6VDJ_VdGg^&I4bG-H
/H)PUD)10K=O>,RFW-#d46M+2:W3H5Y)/][5P-cUV.LMUXIRgdY.4+)DG71[KM,B
[dbf<R3EJ6MLddS9SHGc9We&<_7gJI<WP3OT5)]R;]/@91d6A6V6fDP5cT7BFbcO
eeBMIW8bOFG-I)+=EQ#(@KR-aWVVU7]V\7a\:;4.a^MN9Xg3I#_;,C6Tg?W>NE1E
(Z>+<9.UE[YV)^XcP5_NcaK&e0>1eQQ83ZddEK5bNH3Q:QZ>T9U#_HGWP>1>F_V@
6NP)1C[4P?BX3&JRYc6d[I)N8</78a/K(1)QAII9EG9>1<_JQ<3)ccNWUU8O7?4\
B[0W[Z)C1f.;2(DNR0SB^G&T):bYE]FNOWg>W+/&8a7PA5cI]OaZQgfHf/1-YGKM
\.3gNDI5AVD@T&#6A+C82U:F?b]\Z)CeX,0CCB>9OY,.PJX-IJ\A,\Y_c),D?3M\
C02f-<-X&>Wg[G^[A.gX2-eT)L[GKR:-TO#8.?MZ.RSDM4D_YC#)LZ0]AV<)&)9)
\&\310B1H95F>,1HZ&&R4]R2J>=OS+A]UbdZHG3,V+&Y(7(MgKC5F(8fQ&/??L@H
XPG.()52FY/SZ=Q?-E<(6ERO68FLV?JO;XJfF?<//SLH=b&LfPV]7(@02:,HF+56
5VO;AHSa]MgS2,fIGdTfF&D,W.^)bSS9b=d6fgWT^?d5fTOZ4fIGAWFPP_MJRaF?
?cS1T]-\_I)?#H963FS]E9G0O:91RW;JQ-c;&dgSQ;S<Mc<e0.C=B[G[4J6SCEDE
;<1AINffX:<:2QYb(#6,F=X7;.O:9XM21(D#CL7>Z^S<?ESP0d[VZga[+?Xc=KE)
+eZ-RHCK>=_#,AVE4SBL(D<N;R7D<94VR:VQdW>#93V)>aN-+]^0&f):@UBAG6FH
S&-XJ6\fPcWC63_M]Q-QFa+ZOVFE6Uf,;<FR6Hc&@H\G7;a.LeQ0S5_NO7O\b_/9
,G@eeeHd2N7/^]Fa,,K]F[-8(Vb;f^Rb2OLAef7Wc70NRf^Y1?9e2K727/EV7YMW
=)Mc+3;H>XO\]BA\Q<=S)1RQLO>H>g_G3#;G87W)cDC,[9,Ege=O-bSN6Ce/T15O
?F30^456b5R4MdK)BR4\YK01_&=Z^A(WO(=[b<:>H_e(P6<?dCWY[6GcbY>_6Ob5
Xc52J7,WLf77:JXL<9]2)f(,T>]-@/e@HIbPD]2bJ)\=Ibgf/d.0J(GVd^-O3&L(
g9GF=BTNUP@W>\,Y)GA[&6,QGf+/9[3]VUeNX5NZZ#)O+b1,KeXDN]XT<_&-]&.Q
=LN>4H@N@?UGIa&@?.fUNR-=&WaABMUSgRK5bWY&U94H[AM.[;T467J.;e8Wg_.J
:/_/cNIJ109J#[IQcD&P-M><2AK()XU2C[Uc=_FCMTNJ3<CALQ3Ac\f6PV[PY1=V
H7/O]GTRQ:OG.WP@TO]?98;AYS3G7<^VAJXJ>9RFd)EZAbGPF4bCgQB+Z:b96=]g
g^PXeb?QPTUa(I)bP/IeWALD:LL?AIC,>?5\Q>>6gbfIcAB\\<MF&S31H/acR.J>
#gBZ8Yb0LQ6dW]Ve@b.?]I^dCPc).XKQ3]6V+&HI?WQ86GDfgc^UQ_OLJ+[0Vgag
;;\RIXQ=<XM[B(5(857W=2LGVPY+R:fJ+dH<VKH3[;S@&]#,P_/1=3-FW^YBUNNg
9KgWQ=U<QMe4+2UdCNS8#R4MIb7:3QAbc6M=SOBg&0f)+V[8U+.-(7_B1]D?6?;L
R\PWd=J;c,[B[gALW#GC72A(RB^KUD-E9d;OLV,g0FE]>.1b5;WFcZ-GYAY,]FXg
K]5RM<(FbfdfUd?P:1&Hc2eYd6#2WK1Pc5c1+NI_GN.2WVb6:82P694S(8,4&+K/
J2UB9[&.PMC+MAfa=34F-e)4b32MZeX3g<#(A9Y0:LS/:BgUEK5@VA^)@\\MO^1U
TW=_H\T8E5<ZRKXFLY>4L-g,;Z2EJEf,G?;f^a:#fNTO]A1WNPI#8LL:]AQ;Q1YU
J-@V2.[=/RNN2(9)dQY-.H0:DI+EbT46E/_V#I.Dbg+U=26GgUV3D<^_S_RaSgb,
YQ?O<O&(E_f&G75\MH+Dbb<XB+PJI1[:0Q,9=<Q,M\?QI1dU@K0E;Zg&C5VQE/87
#O+5c2;:W_8Y^@B#937XACT<MX5J&H+aC=HLGeT#]>:g3+VO]Bb&JY;Y8+FR9\VG
d6H\S>TE1W:V][H_L1dX(3TeL-PDQSR6b0MZQTe#6WDQE5,MfR&dUPg#QQ(N>]A]
8OE8H:1B-(V,ed(5D-(UaO+1bD0a7gW@]=BQOG4T>QIWT55T#DYNKgBW[-ZXWW3&
L4:O8R+T,6>\?P.W2[IO-Q,?:C8@R70-B.;/2#HK\g)&MI0U>GKJ6AWd-#^VK+cM
c.O4X_5CSEQ/SUB5)AdcY,2N)eQ?SYM3eJ4^]HTC>,G138.a:^G]bc2O82#?e;PS
L8\=cZBV=>aL^K@5A4#T\X-NW/,ATWFIR_VD##SQ8c+b_.,Y#8.,Sb8D;PXHN^]G
+:d0XOeST1e]TcW\8[EfBZKK3CBf,GgS?YB.P^eBSa7b?=@MW1171dH>=^9@BYgJ
J=:ECM=.?4UD+OUf<WMJYF.QE0A5K9Cc6ag]S?@907P,L)3Y\)C5V5>2Q(8IGNMK
a,J^c=M80I00<QSZ8KCZ=Wf-1F2ZJ1&d2V\/@,b2#=F6C0OQW[N2beAO83UVgWQJ
:1XC7S(2f2_a+Y[O++6S,6EIU9:F>7XSa6=\GbR-))P/Q1E.2YLcO2W[9S;[UAN[
1Y+f,fU&>.[PJGbKcLN,5:S30L=QT=/+<KGg@0EA,-EJ3N(9.d><5K9IXIZGBZRF
e8aJ0L-7-_I;=.)#DMN+Z8<_ZAW1RK3--aJc\2ANYE>H?25Q1\RfS::RXBe=4Z)A
e>Z_S&@e@.b\LKHH[&E4(X2>c\a03eC)29^g(W&P1gQc:P8ee4-6OL@X@BIUK7I5
f@\<RQ#1#W1.>_dZQ=AdD9J.5f]=6:T6PFTEB9N]@B_dbWV,SQ#DLP+?e2LHN##S
b]]UQ.[2)4W@7bN/8Y6PQPX-fT2ZTR\1DWD6SfSGY0#1SJ9Y#)79X9@1N)eTGW;-
AgHYL3T5F0TY;3OT?0e;36=eLa.RGXG-a/2W9EEH/)NV8b//;\&92beLQ;fYKWg_
8f614@6@IJ19W5_MO5]_Qa,ZSJW?dIb22e=&WII3d1/c@WXG(:>Z:6&WJR7)R6+&
BJU4Oc1@QAQE7DAEa-/4RC,]^._dRS\<7<GX5O+CS:f</HX(?G7[8.?[,>_XE.:V
aeJ]R/HXQ/,,W=_c/CC#.CK(;04UO+XeLH3T@d5/.5\_Q9Q=KKXa9(fHggO]<?Tf
1,D3H;I44e7D[OVag5@P;JP@G<WZX,W-gZ;fV,XR+K)C4b7.3?fZ\Y0+fII\.9D8
/?J?eQRP5SE\9[BZFRM\\HFR05#a[UV#SG6?ODUL[6/H,DgZCgO\\=Q+9,2b/e5X
U@>GX17I7B1.d6d<=M8<<0XU.bc:YaLE4FR6+d&V-?_K]][JP/@[Y=<:ZDFS?5&e
^)?U[,VFYW[I]DPU4]O:;9S)c2S;RZ.dLeLUVOWC5)2=KX0_9bWI]YP+P86AZ:GE
T9?^OW&-9.Q@gS(DaF::.A<G_c(V0H\TLJgaG/W5MI4d>e,12)8271C_\2eBgbD7
EGeU?,SS-YAcVHIK2+ef,I0B<XJF.,Da)8XCQK:??U.T:8DdbT,9WB=HO.g?3P3c
.>.T6)J,_^CI4;V/#R>0.HKVT@M[)AP+Waa5WPF.+S.?7:W9BC@V:-gC+(eISK;0
2#LOHM<-V>\\d[KK0A6Z&(gZA5:40g/e/=Wa)N&I12UIPEV)GAgHIQ4N-./S>3(H
S+1U25@2P0V]C82<HM9:8CBaR68#&.=4RdCY(1I7g&)SdgF.;Kf/KHQgJa;_XA3K
8dG1UbQLPd.b.#6MH1)1e=Dd.f<5OPEcG43#HTI2c.Z#dOH:5Dd6bGTIUAXKdRNg
B51B6)eMf^f.;]R?]b@+]bL9M^9M6KDSM)3=b#S?CINU3GV[2;@TIULS6e8B&=:?
,Y]Y@]fH)[SVeR5&1Ka+EeA3]1^PLH<VFb_1Q0VUEfMU[4?=XP_^[;5AfJDVH_W:
NS+#8f+/16JgRW^^&76fR-c76[<V&D2U7dR+^b_FB3S#;4,&KH=3_5R.]F[f=:PB
:5TYU>3Y2AN3#.-FWeggOU)Cc>]XP7,0UE5aKTB,V#?Y^+e>6L;J-?2@7HT#CC(Q
L0MJTY,K1J58IW1@]aDS#/FR?;/0?A5dIK>cE38SNd^_5dfL;COL7.H(<B2Z#(JQ
Ncgb:ZW11#4dA3VR8:,M:;HQ?:@S]R><8d-(YDCZ)):F))6VPV4:I=KPN/85)gQ4
(/g/CV:(A_c5NHI>U,Y>GWe7L=Y#8?b5HL=K4/,,9:aL2X>7=+^dV=AUXBA:[cFF
gPT/7:2\Ue6Ddb+5D(FQW1E6.T\/,G96[-fO:SZae-@A83d82B\Dc18gX\UG&FST
9^T9e(cQSeJNeT#4-VN1b/J[QX1JLVN4&?OWDN#WUNZW&2:Cf]C#X89:0)3P/M@^
[e]6V/H;^IdURHSNDPZ1?-T/8Q&b]?_2]G<MGfP+&9Fd_-ID)Kd.>K[VcMLX](CT
bF^_eP&_\gZ58A1ZB0S@K[JB\f2E.U5Cd3E@Ka+7G1X>eQA?/?+.7Fe_.c2-GDJ@
HT&4DbB>4N^#)e?)Z[_0QT+1^#)d/\>U30DI5&])CP5W#;R4^-2T@&O-:V4?B9EQ
^5^>,\Y@feb+W7+IOI/0UM/W5cBf@f6@Ca5RZM?6D[]L,0MM]JT&04)SE;fBW?1R
?IADF3H9KZOY;#MEec5?J)aW:T;Dc;8fJGfJGCCJBDH57:7_F<O,&H1?@Q>4cZL,
\8g5R;=>S2M[RM#Vb>GG:eC14B+41:LOIU8MI3b_D-GRg\7?;IEOA>D9g\&^JII_
OL_aY)K8e+[_OK+>2=G70R;H@8@LaE7@dD83_?;;B:)0SSa@/7X8Q53=4&UKM(65
Ff1T&08@c3-1GC<G+b=N6=5a?7Ld:U0C?:\6a@U;3KbDBHaH5-U?;KI[</3G+)g1
@XeLcTO<aT_5c#Z5&\[]HS-9b)[aJc5>gU/HEa9^R\Z,.W:OF3gQKMaJ.#<b7_T2
0FG<^c.AK:DHCI[?C>5Ng.MNVWDM)@:QLA>6?Q8e_dDg=F3K14)KT,>6;1c^0D?#
L-&T5J(HI7,ZaNaMPGd0+(5d5_[RH[^^a7&=>/&0fY.;L]<UgOG+U;2XBSJ5P2Wg
_A_.Q\VSGf+W10Z?O=(=P>&Kg5SSegB=BB1=Q0RTV#Pa9)f@+^6R9gQ6?Od)FMB=
.;XM5ff#?S;C&XXF?/G.ZH]-+ZHgARYC[V9Z51Z-58Y6-H+G[MU9OLX?(;KJ?YFA
R7OS[\T&M-<W6W;5X5WNJ40(&\K8JPf)JWG?3g:K#Ec64/IQY^(dfSBH)W(G==\V
b^NQA>.4?JGe8)ede\LX]4]YMHX8R#XE5Z,1F2cHC4G5T]d:O[4)0I4ggc2CII4V
X]Z51N6aVB5PD9e_e(a<Fb(Y/f04S5Q:&:_8MN_@0:0Ib3LMdHH7U1K\eWdD_2IN
IEXS&8c9KW]-E]9[]DE72##]D36J)0,W+));3cb-EO&40L<?J:^Z)ADNHY<.KWTe
+@=L39-\X9GeK@_3G,.[82g;OW=,.G1_fB4=f<fH^>P@ZXWbcKJ:->_:8HG[^+dZ
IQX2DDaeTH#:RUB^+H/XI_5I)Y]?(C,7eaBLV,6/4-&fF11c4@IOJ)@e]@;DY^Q_
#g+9>=@:YC\;O9__8)I>7GXFT^[:5E@GAS1g48C:#\XLJJD3Q7dC<[_R0?e@(gVg
8[[OX_8C38KCAGLGO9?;BI(Z+YLY\F3PM;g+7>Q8+QW#NV:2QefCYe>d,C2\(QB7
[Y09T8=N]Q5?/2)K_I_7eb-Q>4_,<723D]+=_IHE]Q4cIFd;ICP(>UPB&JM6&=1^
#][_T79??;ELa/cLZZ(&,3#X6HCb4W&&H\SbGHF6-N.5^ZLP88)=K4X)V_5fB8K.
E^^>eX>I-55.25NI2130)_KeX@fO].?D&GR(F[<V5)O=KMD2A0;.c[5>1E_/]P4=
AJ^<W,_fQG+S.VZ0;f^OeKYLHfK360,OaA50:2/1@DX1I32&cD0BRO=SLZ]X4)@W
?8)Df.d/@RVe[IGB?NXB&>8C]SLEYFWG>-B6e^48VO3]AQ2&)H]-8D-cL44I[4ed
P-]#a>OdD@:\[L9)d7e@&A1.]<5EUF+67HJcMFfJG;b_J+D]6aNC7QGf6X^HNg#g
5FZfG^Z;)^;SC?);MO+5#Z6U4[cCM_922LKC5TM3C&>g3f-4X+F3,JM7D/QZCJB\
5O&&MD/ZYB;BWOgX?GA#>ZNXRg#g76I#1/1?K2+ZR+PU#NI,-7ab<;)]5G_3gFP)
=Td;>.Bf2BH62YS;KdQaSe@AQ7gJT+N<b<^]NZG9/JF?Zc-6TJQV&_:XV^FK;SJW
)S015@F.Y+b_57UX9=V)[I[KJ@\GMD6(<B;Qg=I4bY0\Q,?S>Q)NJBAIUD0?1I^g
-#X5UE@38>Qe1ggG@39=WGNNN3bJKVD5gNUa=5].47.F,C:^M_3S3\KcO\af?]6W
<KJ4.aBU<=:3F&;5-WZ+JcOXQ5\a]82O&(cZ6C5W?W\/K\7C8OWHc@1L[DT0K7e7
@G.LC7\.J8GEg?Yc&d1)]J()VeS5Hd9[MI2F>UD2QTR(GW8/S6Z=DL84H-=+VXIG
FF(_cG0+[YG1QL-V)SN.R;/<3f=/(_ZA_Re&\0[gY&W525R^B0,[]V8IXAAWL,f;
4K/<,=gRFbPd+HVTFZ&IGg+g.K6&La/0QeX.3WFa-P((I:.fC\,D84PZ\=DPdS1V
g&/YD4Y0[g\^aPBS;Xf&K+O;bb5\PFR2CBb@YRU&R&L+&HUD+;5@]<(?9AH?R<,B
WHF/?Z8H6@SUP4IcFPLX&N4QWYI)2VfOKf<GU47f7T7gc+@#I5-:,DL.-YaL1TMI
,B21U:&DG+>PA3;<N8=OL##FY-)HVeR(K8W+E@c,=73D@b^N+ZD@8/;;]<be_f,_
YLaMeV0Ydc_LTP:81&HcUAfUA>#1N\LYP.W;3b0_[-+-1AJ?X?@gPH0V^IV-+SEJ
I?(P6722ZM\C3O+@UKgd2C45:1B+Z-J#EfcISE4LI.AMJ4g(X)TBd9Z48-c&9]F^
UF<ee5N&[-/b?R-0gAPINgUSJ^BPb^L_?\I0Q47=[fSW\7.RUg.#gQSSA?[,E:5M
Bc/&3PF22gbBX3dgX6-USde.8834#eeN[L;eF8HEbC^YXEeIYI^g,247LXgK]KV>
I5ZO0T(W)=[U=VB?XO;JfNNC72LE];IGfM+U#Rg=X<X;eEH:@9e)(Lg#]WJYWBLf
.FCPX)I36QN3-]g.+&7W@+R-X;3dBT,V9dERCT(BV\X+N9KK:e@F..52R,JBYC]C
/)U]A2(.32ac5B0([6\I^7XL.VFP7CE&H_[/?CeY9[QV_@U#IPRH]U.DE87L>+eA
.T_LHQ=F8N<8.-.](:?A1<TVY@Z>OP?H]E1A?a5e\AX,gF1JS\WfH-@ZfLQeDF>_
Nc+9MWc2H?6T-OYQ75>?[;2K7[OD9N_-7_&7@F9J&\SaEOBU+1e#L29K&3WH.([-
>VDabf+JRONc@V7ZTV8>eH=ZCWG/(VeUSHJ&BeeKV^R@8d)4EH/a;Tf8+=;Adc>P
(^F3NHD#_/,)4]O)&R4cJWaaW&JAAR4f>5(cbX(P67AI32a#6>YE+Y)?JPWMV#D;
Q<e\1;8V^:.FL+:#POW:>EMO\G-[TeXdB[e>?eR#bK9+b.-T5/HXf[g?;=?@e]&S
>8E1TB:A&F]Je[Ue1V?f.X1.:)b##@^<=WW-LM.EaW_Zg;,KOaE9K7E];8;=_@Mc
,ZXC@M:aJ-FJN9I-=V5)3P+7<AD2C+ULaMe2.8U:K807K5B1<Af(^=f9^MWdU<\O
IP5:&.cD#Jb)aIEc/_MY+T,^<d[=/f))IC?CMSgCZPTSY7JMg<GW\6-fJ?OA:]\+
;f?8PEN7f^LGC\e[ggVcL[QWCVR7;44KbMXBDA,2O-;bWF-CV+7,e._O(N8Pb;0O
QBbL>PJ]X^_<C^F66=>fgQ\5)NSLUFGL+4^Fg-(fHG?54GeaJL>C^HZT1B+D<=RK
5?\Z+AQe>^E@X(KeaET:(gYS,HXc+YYX@+IT.]4\ZG?3A^a]O7SFPFM0>:4N)98S
eB,[9KC^UYM2(:c8WEM42KXJB;dg3AaPY+5:N>[7M@>XVBbY>^S>4]De8VXg4&6g
XcUPBTbEQ<GOgRLK2QLKa)O=3O\ABVfDCPg9=\ae:.LXYeYc=Bg@f(0Nb0+@d=44
Q3#&9JcCD=V5c7U-+8.YYb)2f2(-aLa;F\\S&I:ML&c:=X@3L^R?(+YDSQLC_F)+
TX9:63^,DgWC=JdeB-fA>:b;d@U(4I:DL(Z(?:J_Y]Gg=a0=VRWX_ZTJU[,BUCgR
5J5+E0I;Q])35VR(3LfPG#8JJGZ\Ted\AGM-WMPX-&QXfe/UB\?A5P(Z#)_Z),;[
5J@Rb8XE7J^56]Q9P\DH]7#9V8a@V?3?F7Qb@7<TQOO+)5&>LS:PRMI^AWP+F\Rb
:;V3C.M=.EVNQ-+ZWb2MH,b<23+H1XN5&<7A-BUWB>Ae=.^E0FPTO.?5JU@]=JZ>
HUZNaB/+g?;+;D)?R<EY0dfbaAROV+WV9YFW;\&Vcf&^/VHRP7g7(W&)\5(&/Lcc
a@&HD<_B?G3=+&V9fR=#;R--XKe]dD1X_AG/C/.R;.@5C:;](SNS_6/a/cQZ]J[e
:,O3d2\?3gaZM\QR)#P;8Xe\_D_gD+]Ed0Cd#3W>-AB0IE;.X-T3gT6R,=0TW.O0
cY;78\5H]?1TcCZEYI>7^EEb[1Fee>ANgRH^\S)4^OZNddPGbWfZU4-43\<cC?&J
R+4ggE94cEc&@Q<@e2,aF&bS\H<_8>N>A68FP4XNV5D4(E4,[F+/0.KZ1#?G#@42
NG@\Y6/ZL@YYCg&dN3<#JRB(C8T#=N.f?GRgW=71EL6]HV2c)?J2Mc43DP18)da,
g@B+4J7Og+[-KR614+dGPU;;?EQP4;g+-&;_;A)&X)=(aeF9&1D=/=KKgDOP&_R;
R<1,X5IZLCI+VVEFN8Y8GK8g]a?B-P[aY=;K+=1FV#C5MgRa>ScAOI5bd+g=VZEa
c+NLJcD.;A=[g.D9(\QR+]ES/BOfTXRIX10.)B[::9/SD.0-Q.(.[,:E5-U(O?T)
8CH0WQ>@8WO[(RF<1a1aET3,_/-:EaHFEISL(1OXTEE\VC+=:09RY.30BV+V2E.>
cU-ZL+8D/<HDEUL6=>AFWVbgEQAR(F>/>E>D9g=U7YI3UW&6V)7#@/-#]&KQ]fB0
/&?O]f[]2GJ_KRcTfA.MHJ1Y:W6M^L2gBU,O+7.ZE[b1K9cY;U4b.-NXeTf>C++T
UWE[.\</,K>a^/KJZa/5aF[b<b3)41>T0];I\JFA=1(<3=1cJeF]E=01^c-K_\1X
B_=EC.gR9.SedD<BADOD)/I6Oe3N@EK7_6FMLL19(M.BZ2-+F(\RIS&H3>^=:/HW
2V[W6_[-WC^Seff>VN(42>deH5\UV>/AZAdW6\f4W.A(Z+T;4_/WC;=O@cOa29WP
7da+(C=Z^^PH&7S88,^2L55CUQNS9;&3HeI(/PdZ(e<MP;LB&KZ6a<1]QXYT3EE_
g0/R/[<1[+),ONVXbCP@MJ45RNEVb]3:[_F4;d[EVV(2?<DIUafYCJ<W^fI,TO\B
B-bc1:9QE.cR/IfC6HdL]dD9/CJWY[6&a(G#gV0Sf>MMb[WR7_,C+6X>E-I;:_BM
R;R,VH@)L#5A>37U4Zd:SfNVK]@Od,R_Xc9PgAOVIG=7<4(GRP<.EA(49V23(E+\
5=5Y@>;-Fd8W2==#Kf>cG3XY222>9D^3e5/V>R.SNWX/TWDN6/S[QL[?V/g=T(Ue
50IIT0cEF#1)V)2^=CC.Z13d^-a<X:^_B64AIK8e^d5WddKe66SVG-V(PFC@803E
</,WBC2&FC(T8<<-7.R7:\L(N:>KFd?H2+Tg\d+ZZ5IgPA/Y5@^g+6.TGa^DTX=a
A7\#7,6NR[28:BG,9SZZ>4[1TGV7>^R3GUIfAELI+Qb,PeA:S:)J3B>8CR\cE\2W
4KEb;]g7f9+]]:fF.48QGLE(\.4.Z[Ug_9ZS?(d@)BMR6b^AV&&cI=^(,>dOJH7Y
c^12)&;HOac[:KD8/D,(g88@.8f.f0dM7:cH2&2+MJVLI5S^:C#VBeAd0SW)@YI8
XFJ#AL.N^))_\&??^3Z5c2GS9.Y@;1(P9B>e+@6XD,U-=W1NeGH729PPC>FSe]LX
3YDfUL9eC++(^-3EBVY/N0-5Q=YQF55<A;LdZ-\eH];VWD_G_=U(NOZb.@K/[.7+
G7QB)&bMJE@:&Z@=#]OgB=Z&f(&)N<_,):Ca3.U0RNBcbQO?VeWUNCY6@^DG=U1Q
7MOaP8#U-J.d<D-D6_?KA+LLTNLT7OVBO]L=MA]gb\LQa4=;0UKR<g[D#/LK@3?J
/VJLF^Z;2f(17OTLb3;Df1F?71J>bBC+,T1PM&(E/(J9+T2bM[gGDH]UG88(<0gK
<PH3#e,a<NE]X,O55#D&g&Ug>L1;QQ(Q>6c_R.0DDW_Y(G.207>ged4OQb#a[Qf)
Ee5\?[.CWX1+PQHGDP0fB1B+I\8\N]2PNbYO-JA:W]@\HfY=I2dLcH>><AU?EY?Y
;Q=gXX6MA9#GdT=\<Q8(JU_C9ID>.^c:\MQ)H6bF@Ga2:Y<B+)6#8DCQ?_QSWZ32
)IfY1R1e:3\?OQ.#24#3-BW-MLdU>I_ISgCU,I\+YC;&cS->ERK\TO&4(-#daK#e
XLU]LWW&f,0d727Ae-#/I,F[80[ANGT?KZ>G5)N/#aa:\98&+&B\IaPY-:9,#OQN
SH&U\+^eSMXS[T=A(L>U6#HASM]K/J>Z6V4cK6N4;4QcT=EUR&8MG+(f)bgW_B>#
Rg3E&NG<8.X/[+.FMOI=;U;G=e/LRX:We;eY7X)3-,<g_]3QS>cXKd0;Ra_=L--1
]gNJ2Vfbd7DO?YJQD&O5,4XXf5KD\?9;P.(42FH]=ET39@\)ceS;QG)02SK\92(:
1FbW/E_KNV+4(S9YE(MH/6TgLB3PIC.,IB3BZ&-Eca;W1\^eeLXQB)EB=.P#<C[a
BC#TQ?@VSN^d_?N3Z;2d:E0==RdXLZP@L2P5FIbA0cJ&//5=-(GNS^3)&O9_HN8P
bMTdRC.07J?@=G?#,SAb8+Zg5G\C:Z@<)S@1^d@_;7ee4_e:TM[R>/(Rc?=8^1Fa
5dL-eadWRXMW5+9A[YBD.-&>:-Dc4CN<#N<Ab.9;eUGRc3/JbZA/6)Y&YDM](SFY
R0Y8Pb;QOe[E8RA+YFc9+<T2#Odd@g/QIM2PBBFMf68Q3\CObN.H/2f+XZa8)Cd(
KdfI6<.,+T&<Na#+]4W4MMF@Q1+BB9dfM36&FKbD^@@bH]0\WO8FPNS7..I1LDX7
8XRFgFMT3DG2\^D;A1;&BC?,#<[R]+<F)G#J&=dDeVI639P&S5:S(Z+.5<YQU1Z9
&4<28#K;]U7#&)8[QNI7TIU=FR)8-?A55+3/4VEX1U]7WSM]0aOY_RAZ)V-0U5_Q
CdW)_WI5bFgRQGD?<<3/[@495CPUZFAc]]MN4Rg:cM&R0ca@YOBe.YdZT7GMAXaI
GF;e<>fY0SF<=HfZa94IdC-MX]><g(A\Y9UN4BM_^Ub\.9g/HF4F;C-c2Y@?HQ;-
6./]UBbV5,1RZc:R>XbYed+MWO6I0/)J3FXX#XQ7+L]YH5Of?0[cNBI][)1CBVe6
a_J+6Ce:#^JHgg0c-:,#cQc,Pd]<MANOg&bK5F[-VVW;ca8OUC4>?S?bOUQNV57[
EdI>)57.I1/^V/3-Oa=)DTE+6B#(NLc+)<&Q=09F#G?c<#3V0Q)/VYBSc;b;GR,e
YW+ed34F.1Xdd]dEC\?Y26]ZPJc.(f-EcEa7]TRUQ1S,bW)6ae)2WMNfa5\)@3bR
Sge2AMK+Vd)ZEFST>+CBbXYI0bNQEK+:H1]bLTf\D4+QbR;]eW[dF9Ye2Ygg(.VP
@b1_JVU_E1VS?9W7e3KDBcIK:.?[C0@ab3=X3IdD[e4b)@ACN/<AFffg#00+cO,c
0d,1Tc?cE@(]b3L\JBfcA@8Na)79H<?119@&2RO#UgZV9BdNMB;C[PR=,QFE^KbL
gVBb2TGJgg+W#K^-,A&[fD:.(M/dO^)cQ]Zg:?4TV=J\G)[92\#Pb[LUC-&:M/KD
]ba.[9fgd6ZO:OH1<fcV2)6^L6X_BY(3cRPTEGL7;Y;cgZ?Z[=E(8LT/AdRbb6NI
Mc)_HVc4;#bO2NSLX#J_2.0f=)ZEOSce]af>ZZE,DVPE)g<Je+DGeS8L+B:M;]XV
Dg]-LdTC\:5V.+<VF1fWg]=D#9QDEf:QeMX82FLC83_LU-eZ^#7>dd>+T:b+3dGN
E6>c1O;MIMHcET>&+U3NZB7#Gd.<UX\[2P)51b0VfEeHBA_6A0d.Ub;GW?f3WEPA
_M-&.=#B)cB.0\eb,L^/L)I?\]/65]<LCf,5_\ePP[>AW5F1IJ,C/H;S#(9a9LXc
86]:E7FK<7C^Nc6(KY(2[EJ9?e:L::X-<VaV7<>LBe().?)(HH\\GPQNeV/V2G,&
6=J&NFY3(b;A,e=8DI+4T>dd1&<b/Sa/@=_^&,K6&IGD:O6W6aU_>c>VCaf[f-TM
5@d_ceg>V(Ua#9-bRgU_,9&#6RLgN4O+7bVN#9B52?EMJ+5gZZF+<5FG+=#;(Sd)
NM\Ya-O=MQ9PaZIE8G67K6LU)ZEKfbV5ZgIEBI.T9^BJ4ffX),8FWU#0.C^;Wg_9
)]Ic-3&FKOaLX0S0V4T<R6,,Z=V.@IR&)dTYWNd;]RI+VaeUBNDP>DKB;.HS1eQR
Q(b?VS@3cETQ:6=D2G;@,?/@Z&S/P&W@gW9GAWNa5LEZYT7Hc=(DRGIOP[X2Y;62
X7UW&1&IV9(TWWO]27=5F=?L[6]ggUH0E=)G\T_.I]409X&Z6SCXYN8-8.#^75R4
L\/Zf8,^f.Ya/,CC[D5\6^#4AW<F6RBUG#O1_TE#cfVOF4S4bbc:2GZ#2.d]ODcF
Db(Ec8eB(ODF@J/\I#Q,LJBVJP7LVF>_K[EQe1+b-IJ\Qc@1PSEb9g=K+Rf6Z#E<
WSG=P]]Gg5)72TN111f-1UV8[O]3#3E/DV&#1(?&UH:P4G7d094=8^K97W/6(<?=
B.0TO5Kf]eFB=(>XOA;c[gdaVEAbEK_S,C@D/,6NY6H,H)6X6[;\=bYEW\HEGGY?
G)=@+6B/ca.(XebSP#/6DWA><?[V1[>^4QXcW?LDSaOW2=aNU^d7a^Z?d_Zg5:EZ
,F<O8-_cW,]0U/H@APWI:W\&\8;/;+U&H1/WO2^M79WWP)<G@aW#AVT+[U@5Q8R@
fa>6DH9W89XNPOb^4a(0X_bd:[Ke+1TYNMPCXGcXfQULc,8C3f+8+\fULPde(EQ9
S1gX+]N<CCTAO/T0UGHB)GA?064;JK]R+9Mc6AYcW<P_75CMD/Ze;Q=LKI/LN@)6
A0aR>@C=EN=_g8@<].T5TW[EJWX;LTU_O7/TP3/[80NF2)U<XFJFB&2FcKZ_Ob68
6#dZP9H:S\)=0K)bKF5)WHG=NLf:5:)MK2G24G#B0?HGd,+6Vd9Z+Jb+_BA0e228
HdC.d;<39FZ@T/=E;c.AdX>;AIWK3M>a2G,b-5F[W,Z0X8\=I_1JAG#=(VTQXS?[
FDHH@D@<d:@?&?4\;RA:NI=HMc4UcR?D0c\FZFAHd-XL)^0a^KeFFYgWMc9X.Eg/
a=d17VF5BQ3.YeJZCHBJ_>@OV=c:UEGa6NSAf8+OcF429f/3Z@fPJZ5]RdF-g[=X
2Q92KI0bR2+Y@--PD5RK<Cg_#146_GCaaIK([0:_WDC>/CN2/Rad7a/NUb<@F(Ia
XA6e7,OH>YQ8Uc[EI_gPgG(@@J32)7_5OJ<>d,/c/eOeDf_(<+eR=J0[<YU76E]9
O]P0,+7^6e.UAD281SE&XGg:J=faV9F/EZG9GeaT.L<Y307GA&UH8^S5^Hf<31MX
<&#<S_@6Ab9,LPSFX7HZ,>M\]AH_XNC9SH5+(_MEd.:1FfcBFZPdb3\&9?3XOg)e
WEV7K0DOR^()1fP<OA^UR4A7CRKK/Z]PA,H?U1=XD?aRM[.ZC4D&\fN85QE_>2N5
M(:GbFWV-HO63ZS>&E&gfIO4MY;&OGP9g#3:]?;)f]Df]D]4@&@6c09V;W.=A=L^
/\)[]+#>N[2eX2ZUgU_LS+F;f:B6_2D/F7->ee[W:cN]0,M:UB\S]?fLXb)0_IE1
E->K^Sc=\M0cCbR:)X:W1+NO&WO@eI5Sb#V;_QTQb3aRaVL4;[Sb)F0R8^<.L_,-
7D)23:DDG#@\^Ac>/84MOWcC>P??D_0\eNE_f[7Jb:O;ZWR;150F(HV9E3O;0W;Y
A:eAeP=X[G=B88aA?R,?R-C+XLMOP;>>U\VAS,JR^@P[D(.A,c\e#/eSYYHNZMEP
,[XBZN03\fDR-ALUE9G4-[E?&#9d_HN(SeU6<LafCLE^HNC(8fOa0^dBKf5@SB.E
dg)TS9dJMaUbMV=.S;4f@JBD64d#5Q<CE0&d6XO[)DZ,O/7F6cN[&6-Z:g2(,8f7
:4HH-92_ceXBd?d>,BA(1D9=^]W)^Fc)V;N\5Lb>I)W21O;4e5D2:OK/Xa-ScP:M
_./e/c@CW:Y7&I1fTY>TB<^Of6=f3L#,ZN[TS^W7.f142&<S(O9;9O.#Cg^&L3c#
I+8UKAV-8+E8cQd#GEIDF)(+R>/b9SHBP=;5SDG6MeG;@HNT;J]P4L<Tf)E/;H^5
aN.6+eVT.XK:FB,;CcS4I/ef82N2dWcSYUfef>ZSa=/W\Ae_EP,L-D:Y^\4JWS]6
BbX6a<NK3CJ3-UaK2NVF\]0CfGcCW=6;a3eFT?JL5GbJVI80KI+X[gY>1Kb0cX^K
>4RC]>dX)..^&7a,RL-E3#g3ZcJ<;OZ^EE]E3MYBX&MD42B9TE>VC#[D6CDf8S</
4/R-:,<#P;+=I+9KPA+.X1)e4cE7]YO#JG;D)86c/R]U;,\d#;H)E,Vd(LQg9VSe
^NVU>-K;YaRI7X6CJ0U7E:cLTA[EJ/0fWI(/KEXC6N(>5V;<Ad376)9@&KQbc<NY
WR:&3g3b?:NPgW1]eefeO0YAf_<+[34PSTeD[>MLP5f99S?Q0dNQCP;IWJ7;T,G6
fV<AXBG8RIJ=KNE<6K;T?#9N50):cW8VQY(0O)H.TL.O>(Aa90MJ_9]+NJ<5TMXf
4,=>V\?\cZ,0=<[&<O(8gEF5-:E@aOec64,d?L=M5d/ZOfC+RCT880[>&P&9ZN0b
YeCBEGNLU9KE:C8FDCKW^W<>[8Q^;OD-E<U;IR]Dee.]1Cg:35R8R:)8RC^cDHRF
3eUGR2@9dOK(+.3A&AD-]589^EgReNNGLKMS5>24V)GR8Y0F8#<LA2M,4Z4@a,R3
H=UYZ\9FPW6GLMaV_0@D-#E?,#F:E;DPZCbe)N&c1Gf0GLG@ERa6-R:1@Ee\NBRI
9Y+<>4Z,;WCP7Z&/1@<b,N8,a6T84J-GMG>+C,ZD\[>D+E1ZV<VNTK=Caf]?G)1<
=U\/JU,+ZV,)aL;X[23?5J/eQ7T#CA8V,I7b3c/7TTTQeEIQ9BN.(>0:g;f6SDFZ
XSfJ;2JD<-S)?REWDSf&#EAYO0bW4:EG,[;LS.R]eEY12Y;B,-#J,GD()WYKVF:H
5J7_=R3f25I/VCV>b89_C@:3[.Q_&_PA3(>dR8<&JaCPd_RXW6=C\Lc\c:@RRPZU
T9P:)@F1^f#PcVZQI??QUST/aR^^[YBc7[.+WfEfIE)4HK[&W-fY#&;S5I[5eP[B
:R9bQJaTQcA&PE;D,Obe<=Y33B;X9P8daH\Y;7FdW?O:eZGIS>fc,?/F(-bKb4K3
N36[B/TH4@<KY3RPCb6,R0Y/O3c>ZJ-<))_/^T^cbP@K[f,IHRI@;6fZO4Z<L_38
2>IMg:J8BXg;H]c-3dVZA\5GLM3O-bSVXQb/_[ROX,B+;D+3MT-aM\N2V&:?:#G]
DXCdM(_e.TE55U9g1IKS&WbVSb0X=Y2^O,PfKQ3H<CH3Ea-b+YU(dS557d[#P_I8
d,6FVV[WM6aHD6aBaEMDH\\71W@d4HEI>3IM/I/4V=]gR5-3[+Q;?J2G4Y\X>(,g
<Y=a0HbDFU3<,-G9#Ig#CS]/JN8\-Y3@WCFBY>1@L<+K[b86=>C#b3]<P:V4);B?
1D?&@a\FN)=.;FUJ_ICS&/Q-UKY4YVCGd>5JTc^8]7g^5;<SUZK7H[_349:cX#[A
.(&f(K(#)@#T^bKWE;W^Z-d6NT_<S@ZCY5b?TBeHY;KdcON-K+G&M\fQYHI(K.>Z
M3H<a&9@Y3BUJgAXCU</A7Y#DY,/2Y/>N9BY=fR^0VJPZS&<S(<dM/&O&,)+<6JR
?[#N9,P7Q#,5?&>YZ-TE72(caE?\B14Y5E<.(.@#2a3#KK@SNdER#H#f\VB9P8Z(
T&E,;Q12W>PXLf;I&NWH[e0LMC#7fU7>2=B[,3??3SHR,N=(WW-;bO3^0SYZ;7T+
,0=:>&cE)eeV+4&OJfTcKb,4++A72<<ASHE23D:ZI.O^ST&30XFC_]#a+<;;)f)G
RCD,bY[6bW&)Y3db>&K?:^1QSO:/:3N.VZQR&f9]+=+C2b3f)g>646fdJ@._BO.R
;PIH-LB\,T/9A?7&XE=YUJOa.(MUP=Q6/KMC_K949\R7ZG.T)I2,@Rc-;<0DU7/d
DUa^6Z=aI<a6.<,>dKa9\D6XZBQ0bNL\2IWA@GZg9_#[ZJAKTd0;O^6U-eVgIZ(W
a_VK/8V/)HfK>IBM@R8K]>,N_?J(JQXT>BY>62cOgJ-XOX(,660JcNPG)@LXGTAI
QRMUe8SI9&8[gHf?K(E3=.fH=&D6T_-=0AaHHO=9_UTB::J2-IH=BZ9S2LTYX?92
C9.HG3:E?OR:NO2:H8T0CS2J9VC,AC&T=S_e&cYLJJF@J+dZ:E6b@LeeITB_QbZ^
DCFJCHf?YO3RGHB^dR/_\H;[E--O+]&bK(T\d,JG^aXcTW)_QG<4;9@ME]fSfUOC
YUS[9?KZ_.#3\&D7B\cS.g6>N033FfCX,V)M.[3>e/=?Z,?g3,3aEYb,=RY&/b@2
P;\[Pg:dFC@<XB\d@U\W:QdYI:P>X=8/_>;=RPXZLNJ);&)))dLeX,-K>UI5ZG@=
8Z#/AbX;.c]0U3Q1;S5fMGT^9U=GD=\eb9&&QZgJPc),K>=9E)AV_Y/]JaTBbe6D
Td<U@O,;7+7fO0g,?YR71/^&S)SCf7=@;<a=:4>?SFRZ+)R+?2cR;X,H:<9J^B8d
0;OCU1eZQE;ea\/a-6ZK88_ON>+ePEIW_\I9BfD#J+K/,>N[.gOae9J/9#>N:1=g
:111F/2C=5)XO/;L61U2-\\G<SK<^W4Eb-[X]BTC]##1>VE8JYA19eY^Z8\#CWeQ
6>#,=?d&aT.XIfCLPOF-UU/dZYOA6YVXG;W9F;S3.#XS??Q(SP:2J2#N@;2LS+IL
HP^JSNVP[gE_/6/X08eO)W<PTE57<R5:cc[=LbXUMAJ6Z/K/HDVaQ5;.eIf^J-gK
::15E7AC,Y[/9H6ZW?3.4F)A6O2G^HC2RcAT[RK;&>>F]aYZ<3YW@I\b6eG+>V[S
/2fKMK6:O^_JI>b>?<H:&IOVe>13X(,U3,BR7-E\4XXY\F52\^gUEW,D7YLdX&IY
^f;edeRg]L;5O+[3-+^a7TL\>fFeE]3H-DW?5d3A[/,2M6AIL+VdTE^1\O&gFeGM
+;9\/<ZAa3Ub_H^):[\2[?F_D3X;6;NP9Fg5[f4ZWQXHM/ZD;Q<FEcTFF&K+V90-
7MNNVNWISeBT<2c0]/4-M(aLY0bP8;1F3Zd]BB=/[F,f[_CeX[YHESBC:c9T.[84
Z#HYMXS8TePdF^2W3JdXa6Z,Rd]ON\?^SY=feaH_(EcA78GB2/\/>)WgKAYCM#=\
XMO9#9^_gZZ-VE20YN6Pd,g;3?-M#XdVJOeK-4)e<Z+)f3V\0H>EL@4OIG3G/Fb9
HJ7FgX4;?/VWLf2G1(1Ba-0c(:\/C=7]&^DV&,3;g,XY^)QddDDaCJ4ST8eRE.TB
:=Z2Bc6&15T4>2C5HU.FWC@X@d<=)d/>?J3FI@S0f[4]cG2Bg@-.XKYb<0U\3_bD
g-9/SeU[ER&d(-GMFF.88A>-ZbW>e^/e1O+UT\M5)3,_)N#,f&^+?F&2.3dI?c8F
0AO(D0Ec?EAIfSB:5#2<BER5^9W^N/VH>P7f4gEb;:d&75VV=dT+^XW\^DVM<S4c
^4/3JT5DU3L.43P2>C\UbOP/#JVf74gA-[LGWZ1X?B][dJabY]K?7I?ZJ?8#SC+J
6ZMXc2D6FM7K4X=gSK(:UQH)Cc_P^A(]Z>K5:f10\;=N#_4)WHgPd\0KE2-V-/7B
XLK#<:FN=a_^Z[O(EN4.a.IXUaNeT7CfGP<.KYe>?T\1+Cd)_XGX0]@fc7K(eg;6
.aW51W36H:X4Bb8?XCg)?W.C<J_YU:cAPN2FZgM6PHaT?D2[KN23H=906R@+0#]0
(H1KL#gaf?aX5YH.g87Pb)?Ad38AKPCVcJ9(9(;/:U\RGeQJDBV33B8?aCJ[1JWW
cSaTRC0EZE0@]V(.a<aRZaG,b1SbRL+cg;>,Y/SP^-RHHLYNNbO(Z3OR)Rd:B^OC
,#e>16AU[+0\S<GGDX-H>bSR8]M)\g>+BUe+;PDg\Qga8H(@B2;1(IO1d.&GWI.a
/94]G(d(9.eUBUJ+08Z^YB78GXTEK<-5++5<;(&/3KT_X.],7eE\.]1TgQJ-SBd)
WXFAVf#D.1J^>?F4GLT8OHTOaMKKX^(KcgBEM?OH:^Mb&J#810W7^]>^>?:L9/(1
aN4NAA(b?UVU\G@K46Qd9[_dWE&H3)bd8DWE_VJ9@Mc<IQ>)1^U1IO8_PP#>=2YC
R7TAF.Rc\b2\,9>V4X&/c0a2^5K\TOBU]B]#W6DPWPLTZ#FH9X_HXI<Vb8F\4K?c
6J).>&PV=9>JWY(^\DJ6X,1,+V/K9/9T+8d_3XN-e-R>Afa?G,Y>AB#S8?2L2SbI
e,,13-@1+^I];D5fQd<:OgF@FDCH.(A.KH@,He<.f5/:C]TWVAa.OOe/:-e[YEVT
bT^7@>_)M48^,KRN]Y_[dLfd\W)7g(.cXOVBN5+#=f:;d5MJZ3S(6GEVQ;R(Y#(&
[H7e>DBD;J<J(Z_S5b<))K4B9TU5CI92==6^W4@8HSTAK^SVbJOX6SHW(W_Acb_:
-58\Y?XL]_K&Md)gO3VW,G=U>deA4T,EVS#13PH^3;H[5Ec#699b9,I>>.?dEM_T
5MdPLTZ_R>#c_ZZ7K0N-6UY&S^/2XfAB]J#JAIg\XV;9d>9]Y^41N-efX6:6GOG,
<,Z8e9+e+8EG5cOaHVEc[.YUI>71GX8EfE+A4.fGe]/Bf-&UK:[VV/dFH5L9]eP]
U&-Fb-[?F=]++WT-FA0R;O4C)#5)4bA>?-dbd;]IGGKK4><eDc4gb=X??5(c7LJC
;83HN=:9Tc[(/ARbG=7bgA.4M41@3BH1Za\++N[7[?)QW\#6^6#Z(=dOOP/Q2L^B
FH<-O0X].cV9@<AJC3E?ENXEK:^[I+^LWOF6K=C(I,B#;^WL)LOeGFd[-#;,#?BL
9UbQUV?eC1A_,cNY&Fe26R4g.=6N?+Ib0d_7NLP(ZK/#=gNG]KD74,W>c18>>1RZ
DLR(G^a-#2>V3)]gd<ORbU3:fQScU]FFOIOX<cGFRPaW;[<,#[TI@=-W[>6LTHUd
3Z6/T16LF_TU3cAY:ZbK3FKIV<URed:L>MAg>L&IaV/1UQ#D];SH;K4HB2:8C5D>
V&\[EBHG2Ve5>4ce_DB#&[R9K8;9R.c4dUJ\fIAAR-[(gTQ@bC0/,Y;6DY^3VT/K
QTR7YCZ.a4L-4?8B^Y-O(7KDA(0;eGVK368^0-U96eF2b@1>7R[U^(N3&:2[2dK2
TgP8BN^#1QAO:6ZYKR8ZJ1[V]gd7Y[_7[H;(+RTV<[5abMRD=;I_G39(0.HTWTZ(
V/;/Ra9,_+<>?6,+d.]aDM^V;5g4^::AAR5V=c]2\JY3NJG5I=]8WM&-a:1&NfF;
L/\#CN,[>X8SGAVL6Y\7gSTNK;G3<;dQJ7>Q:.E7P+<JfSd7GO(EB&+>XBaP2d\S
/6cNQYb5D6S&GD49D5/+6NVX=46[MGG<ELJ3-AONY:OW?7E138<Ffe,@;\T5/Q;G
;N_Q:9W9a#F.EAcR7Y23AOAS7TT6C[&1>-,)[A;P9,g_0QS1T=E757]UGL50532G
VT/U@a^DTF]-LVFB<D(.:5gg-F.FH(ARZ?KZSSDR4V\5#IDYJUb@4PE1Vd:N1;fU
6e(-[4I_@+B_>.UF+ZU2]G>W,aMBA\648L-K7/f-3<7XKKCG^W.IS.,be+.X^2A(
dV?3Rc=#3b[cBEB[g[:K&EZ1CYdD0F<U0PK4EPD#L0RLeYaa+\<-2(I+=4630/Q=
b^6YSfB6/OMfTdeD[79+PK6V2J^[e.U71d8_HKNcXfE0D6D<&3>N[C9D[L:7TYAL
JEFR25CWN8c^:7[;G@F#,.ISa:(B9c,=6^(OA4D?,.](R+#(G6^K.:8+Y91M^2@O
gc<V#^aM3^4MI#V1a@PXXI3-ZF+#3&AUFaV\OQ/&451g4F_faB]AVL/GTH)J.8<:
79fB-MAQLf+9G4]Z@8]L,F<3&c8g1_;[E@CV^RYQZL#[0f0GeI7JWASg_b4).\)B
QJ2?\T@dPW.J<>H1LgeL5WW]0-N:PC>M&8@&PeKI.cL+IVf<NFdV>\g7]RD]?0-:
QC2c,bV)0JFJD[(.Uc#)O3_JdR4d2#MIIGLGK1<0T#X-cOPOJHIKe=Z;?,CU?RBb
_Y1&9C5C9aF_+0QU@bbfQ[?d<E_-I&N7T-JTG.]JCDPF(R&@&MW0Y<@,UH_(J0[K
#D3VOg,NOSYa4BFR:9CaYbWQV6?^L)H#R-47]YEP;TQE_2,-.CG^X#K[VPa,@PQE
_#]EBRVYABG.[P=P7\PWZ&f1M9c5.ONLFZ31T[?LX)d/.53YRBE<7&0cUPTO)[8S
1M-EB,MB9\;7.eWRK(_&.g32J.eI6bNG:DP2I;FfE4KD^O2.dcA6G\JgU(gA9A(S
(#_AYBDC;T(;AK.;;f340J2KP(O;S^^;\(KS:#^/P0:1?MU?N@^?@+9#Z@ET3Vd#
eD(?97QEaB+D<QU,W;-58f1E,@=RQLd@M[G+F/7^Nd=Lg4aPJ5V3KW\=ZKe+c]G7
JFbVCN.-JISNMJV820PC@EBa6Cb31150@X[6fCBdJS^O4@[D_]K&Ke28+G^/V(2N
KcM?._TW,Z8_<F(YUP1@VP1&J1H;O&Tf:U89&G+Z+;cId2)0<:8[de,9,BW>fc;.
cRBEJZ8^IRc4^NDECASL.9W#4>dN28IDN6e<#F3S0E+HDZ5?D+\=J:#=<TL#?JG9
C5ZcU,]3[1G,8=;.A;D9E..&@V(E_.A18X9L4PWA/BeYCf:FN.b>#La0QR<AS5ZH
1)913dN8;O)EcS\D^bE,d8D:5@8[#H;]FT/(\7\2\U4beD_/eLM[f2#/(PD8BV,M
FS\-]OeQ.K5R:;DH+acH>=^5>=HSBXW#QV@G)\g_[&U[DXcEc)D/(fRTSbcT@\[8
S,SPIcFC5S2H.JY[ERU?QPaf;g>gRU]39^H3RD(D5I=(fT>AS1gS5TLQV\?R4VQN
C3P)8:G-D[fZ7U;0<Tb606-f^DD;O4;]HE>[g;7V-&/G,Od4M<Ze,3G44#DMQMHb
)D;+9C-Q>2=+PeVb;8O+?ZUIYOdHZZ0CgIOZV47,Y.N/+R\,4CZ/dWg-MP<_4?Y7
/g4S0gO+6#V=DY<^aaE<[-MU4A3-,2g6-bdFBBa84T4d7a):/XYa;ICOY9a^)W;S
VWZgBRS#2+;+d-ZRcWa9:8<4ZAN]?R,_[V=#L[0K)_\VaN)J#K4,]9S83-eb;9I0
+\UbTf#K48_7f@Z>J&g[L^O0J+V8):aQa83VHLa?KUBdU5RR4/2[>2b9a?Y2S(Se
6#E&TI>OTI9S]fT?H2f&\#KHN;ecB9c=V9KCO4g>PK_,9NK=XVL&77d-K(afKb5J
CEgeS)2)@=ISMf].f]a[]LS9NS,4WVRQ)_BTJ=VFc-XF;O2F1gG7I&5c;&T__fH<
f&D2Z7fd5W\S=>L,ES2Ha7YPVa8aLB7_/#286.90#EKW?#N<?YN)QSD@=+-B3?/&
(\A_Ne4HS(D#ZTH9d&6b>&P0B70NSfcY#,K9&Q+Q_<L#X/KG9_U8@SFR4MW18IZH
PFH_55d>L.K0cLS+OFLG@9\Ug&&F7>ETV1EVc\HI@FTA.3-FCU6-)cRD.V8X:>-&
+b^BV[dADCId@VP+g@6,^,JIRL(5CH-_6=e^B@S/=QY4S5VR/]R0Gg#;\&HJ3)dO
U@YT4eU(K)e)/#[U>._25-Dg^cN_L@+)XAEZ8-HbW2)Sc-a#Y_=Y)IYR9-R2/MB&
[FV9(-JL&]K942D3APSf92>2bG3?ZeAQ[+>L;Y&I5+3^E2^N^.d_UJJfM5f0^RO0
c15175QVVKO0cLDGN5[VCZ-+^/c+d=gaM5RH@[=<gD<Q;MBAFJWL;#gdA6)TM-De
S&5FY2XM+E<f-SB5+N.E6R.9BaJRQOT?T5W/U:B1?KW5bC[U9\7a\T6UTG^#L[X5
?R</.[&)B?7e\0=#R>)1Ng2LE)cb44MV._ZMETN<UFf0R>@.<?A.X#LT]bPMPb:7
8c,,->B8P1@/#:UZN[M:5>O,[Z/TNCE-X,)I^_d#9)A]e7JO^UaeI<[K:fMXK4+7
Nc+IVJJ0/?a9eHHX5O0XbFKeCD<\L@[\W)]G6.EUL8dV^0H&8eB,;L5C(=[^L#Ca
[Y-;GIGE(@:5],2D5LScfYZ1+Tf2.,(cF-GSbbG<D=>DQ9Q#ZYEZH>&(T-Z:]7+2
<@-[d<H<1Oe6DR\g0-K9>&aN.5_BE@G2-b+cD6AN/>&J1d)&(=cTP26UKdF&EAV=
VM2(5DUFDefWaMA_P-(U35AI#0S.(5N6,&O>M&ADPB2;9g^/3b+>Y/RcD,.;W-UZ
g?ED9WVa&=Ud/.-eSD_J.^&M1J>VN79dR_YE&c#Ub+>AKWS-LU1P.P9^TdV=39BF
M,b[&<I&^@?89T>S,baA^c\7eNS-+E2O-H935^,UWJ;S#UQO[<W+[=ag)29#>#-N
(JC@=/dT[H\\@#:bAXW[I#2,]QE03FWg+B>Y0ceCF1>5a_>78D[@>D_<2\N,=8JX
eY(2>[GX@2_2#A;G2DP-A7_8MKD(YDfG;ceK6^:RV2RY_3J)ITR/Y#fB^6E+5^Q)
F.<9H0VSY_7\9NIVQ9-;CbFUT1A<LKdLZ:QU>_cE;ED1dH16DUSSK+VH34<Q?SdG
M/K,=G>;S-KG]P86V-\3D4LbdNUVbE]JZV8\KT>9]gCd8)/P22/[EJ]eV[b?DbGZ
eHd,6QR+c(PO^5:?X2C.2d:,78H=)WH^?HHL6c4#9DGB<J0B4c1fRd[I:&<NWNZ[
+Z0EFI>c^MS?S@Mec(TJK&OLgHdC?&FK<D,@cG-IW3N1?^T\LV;L=Q<b[3/<9F6[
\a/(;1U(Q8DS&3Xc+@Q:GF?B_aJ-6a?V1,^-CR6SI(gIUeE]a3B\#TWd>3LUVS]:
6]9U@BSHM+IV\cb13./dK/.EH&&SB:\EB969GZ<I]NZQM.T#_@VHA)0b#_PSebC&
E3B-LUNc52[SY+BgUWE5^1(F)GY.+ZF#I=<X([(O-OI\WXT>M^U_UfAV9?C##cJ@
H,dUH9CP:a:+H7T/8cP&gg=6fS[+c:e/7W#b9?E5I(X0(ZNS@GVQd,D]A-J_+38F
ee0.&@3158aNU?7>79(W>0HV6fD)K.1Q<,I.W(_F6cY#5E)OAXYQ[S\M94L5+<<E
,)SO.F:.SL+@+]]MI9Z9#/OY?DOd3K3#e^)BKd;^[dRTF@]SCX&aa/]]EFSZE&<^
S/PBO.&TR8G82e3/&1[HY6<T>[WNZ4<WWX=:/[VYUMYG]N,UbD0[<.2@)2(0AB&)
)00/JfB&PdV(3K9P;Q1A;c0R>4P8CWYcL,1[BbRG]/WR6]65V>c\TK>,c:D=g:89
4>GE<De-8QN1cXE7-B&4IJ/[[fFO/USZ]1<aGGSJeN0A,H_#@O3)&EB1GPE0UFc3
/=HV;>+PfF7Hd1QFMM8)a/43A.<]N)K.[8=9V[#>?:AJ+NZO?dU=5>XDRX2&bcd8
d1?9ca[73GJ/Mf^;ZDdXX1;2AB1^>6,F((9#c/bN;/>D5>9@4F=N54I-J6+)cFT@
K^8I6A9\_Y6(T4KFEb>0fX,MS3.<,IV\5-W:d30;H#MbJ]9N0PL6QbQKQ55YcVI(
&N2XUD@]FCeIBULK3CMN@,?5BHNb97T1]BXFRQ.e.63aVDT4Wa<&UdPf#)2PTA_F
^SW;d&Q@JH[G>3NQ191U=fV4[GRg4:Y/9+2&34SJ+#.a0SeG=0D>_XIfS_5eQ.Sg
V:WV@2Z7;R8bG-UWD8BFeH,aI512\^/3bJB4GY7HXaX0-H^aPS6LD)^&>b2B9TIa
U)LCZ_[bQL?fdN)A2d2><1I/(6[?aJ=E8M,;,<0)YBNB3)II=])O)U4USY#8<0G;
@E;A@7Z9>5,bC?3S02aU85Y;@bdMTZeQ17&SeIY/D??W(:TSbOY7W_aH>V([VFIG
(9JVZM-?[GF8?\_1P47#D80(@=QJD;SED=Re8Acef+1CSS=9,D&IV97X_\G91AQ;
J:bS75=4J<EBHAfGgXb3/9QcTa:BN3G(6GR8:V8(]8eOS^O3ZS7eTM8_XVEb_L+D
8T7O/TE;fGS3HI>PCRbNQ\S4PWI#N:97ZQ_E.N0dFQ8aPNV+5749\2_V^cRT;7g/
V8;^XdHNA4:>cA5)AZV^L:&d<G7HN1)H6F3OX=F.NN2?=;,@BVN1^O5FFcZ8+Z3M
EAUBMAQ#C>2eSP<YO?d2A/Q@H/5QeP_M=J^)Q?\TbLXPIe/6SFMgU,50)Z8ET<D<
(TZ/6PV+<)<6WIe;8bB@:E2Q7YJR,B4&HI2P]d]DPDD[E_g^g1\.]-,-9/DEFBD1
I]R_:9(\1DD_D@VZ@AZK]gPQ5Q+65E=97NY/\0G7@A6?CYg]E]_KRZDV7?3X/K]W
YE_cE(YZ1&JVe?c.E[DVE^(Q^.#7QIT64aOA&TdQYIT>,K<8G<#U-<f1^@#e\-e-
<AGT@5[+9(4ebL:(51gK+[0.B91g@L/C5]F)&5?:[7?X+KTfJTRFW@:U468Q@Fa]
cLfaT9@VXEXD?X3Z0+Y-CA[Rc@/ND9V2B_Rc&IYfC=STT6K79?NVF-MHFO/P#Be@
JT_?:D6?DYKTL>5]L8LZg#S3_g0NWb9dga2S0Pg2ELf^?42SbHZ=A?I23N6N>9Rf
M@&JJF(=(b8EJG9c/V@LcI8@+8f9X#MK-]E9g,4)XL0A^0H^>T_\W]a>V5cA,=>2
LQ16PHE+<7SbNf;_4R-(APcAL3RQe3_2FZOHO>2P)+DPc2d9@bHbONI[d[R?/LP>
:[EOQF^W=W?e\g[X)&eG-,6YCa08aB/[9,6BDf=;aE_.HMH\8=+V-@R]O,?BV352
Tg,=6HY3TQJJ0)[MBL_d@#Q]VfI,0.b,fLg<U>6Ye9O0ALAM6g[<ZX^PWd>ROXFH
IM/WDGCW8F7+I=C8^F_eJAcR:RJ9L)cA\?U^83&7>&JO,GJ6H7-P+&K[ZO4-8P1/
YIS:24a#I4ad;@66_2^#b?eM(V[Z&A#/#/Z8H,M5Z9(SVTCUgNSgaOA?3J,T[^T\
?+X8B,7J_]80cSE(L51gLMN:ROTJAW]5)W0dEG/=a3K)&0T)])CDa)=JNUSYAJe\
g_BIW6M9.P0eW/)05)?&TNBX3fFM;H@FU/3e;3GUC/6a^;fHcdQ._PP#C^T00DME
\HPNK&H5+&=7GdQN+JXODF42.PF:0gW[Ib-3Q^g6K+:(MF>GZ4PD?0Q.[Ng_?&I7
@U2PSZ[KH8X[G_-UZLbUJY0TE7cK<Z_<@SF>_TFR]Nb]dc[4M7^b[D-G,5g.cN(a
M8b?XQ(SD^VM5D.8M[RKR(BP:L<8FMXMUQ/8X,1(\cC9E4]@UP?Z7@GPQdD/cJNN
[cV6cA&O(@L@S?WC>&QUdd>TU-BFZW3S1.^X22\UF^@Z:2Eb8P?2-7)P#DUX=#J4
3J+MBX2^P3#]-.VCSPeENb?dSFFBM)/D>&RD)BaI955\.eB+B5=+23f?K7OXUH0d
PO-8B+(INaT;FC<82_<@Z^A4bf2aQT:P;eUKae9O1<QZ94cgZ;O,Z(#NMgDURbD]
OW54e92XZKA5H^2R=^8X(,L;@JAS_JQ=;WWG@c]NQ(&WBF\W2L,e[&cGaVFYH3bg
DJ7UFA8)Xe^E@:gMY^@]B0VA7[?19^8TgIG8,>@/?cGK_Cg+eDHKgNY]42]CAH;[
7W.eFEJY]?6af8&PTbE:G;c=?91JOf?=8WAF\)Qf4gAE?(3JD<Ye\8189WWEdJO_
0[c1dU71]35-Q4+5]]92GYUQ3^dU(JLSMK/&J@UdQ.;335D;@/H\?^b^L/K[4K=R
95e9O(JJ6J_K@]64B(^CSG6-cK@a#?C^,J>@D5[1O/3bGJL+PE1PS86;gc#DE.\Q
0V^<:3;=&@-Q>X>+YJ3Ce#5,eaC/[-]?bS)<W23^M;A6B6Q.)BL,1_g^O)=6Lb@b
&+5e,7PEQ;T2BUM-7[[2Z^/T(@W,2,6PE8HMgC96_e8UY(2XIV+>W?P)N@R(CJIT
[97BBe/K@5[B.a@EOBaW^7(0KW#g6VATYV#fI_[1UcTC,3RVNC)QV+ZBGI0Ab/^H
Rc-.7:6eYNdI:RbHRK#A9&YD]9JXK\I[bY6SO1?Q>QcUOP.,J_7-GSOP_<)[76eF
KN,CRaggTbDbb1=W)_(BY7Q23N+[&9O?+^A#@0fUQbH^G_f>QW9#BY8A+H./E0)+
K,RW>U=XY+EMII_2\Kb2B2TZ_M(M8K(N?=N\/FUWATCD1.7S?:#B>W;>eRGT<]YX
?_0&\f64_^?IT\=,L\b)3?;NP9V@M4DaY74aNF<&E0+c&[d<O_>_E8K-BP:>CXKM
;MM.].&FcR1LWKa<J?U[\c#@S^IbERFEYBaX#/.:c>D-AeN:/L[<aVT:]c]f>[@b
L414#d<[.NWV\U[<?H^9D/cIYf;MD/+WMZP]-QGLS/E(0BZU&^L5^MQ@O)1IcX)C
0Pa<BL_A(ZX#g-d7e<@bOb1Aa)KKAXR2\1CA8T\:d,#/6V\Z@<^A2#TQG\YQUc_6
2C)GBe,CCZ/Qg9/f[NdOEfG8W.^MT]P/7GI\9:42GQWb4[YVE=N-K(?_73B&E;Q8
D5HKAZKc,7()?TYDG9VV-.TJd_A044E><84Fe^TH^W<eca?SSKR^PNb)W1TcNE=1
GdU-B(?Q88Uc(/?Tg,<G9#N>Gea8EH)W@bVJO[7R\c/a)Cab?c])\Y1A@5?e(e)e
//G-;C,cY+1U]C,bXg-7d&OegV@)Tga-\4NZd;9REfGF[.1(??JC5=XdZ=]DM\I[
9F#+^VdQSK-U+]ASI[QaA^H[R;^PZf9W<R1&Bg7TN@Y<Y:#&K^[GaXNTYJ^#8_AP
SbJXbSW7:Y?Rd\gKCa93D1GG4MUgG;3DR-C@Pa:?#L&g/CJE]fZ=I-5cBdc(-78D
S(A>\,SO8Hd3A2D[K2PZ=JI<,6bgQ4Xdg?./e7JB]U+b<,;))L5D_cJ&H7LEM>Ra
OMCDU58d\\(Md_Z\ZM,bOB[T5f?#31g8CM:2]UZL/M.DJ=Ag)eJ.]K(QIg:T6c5G
8_W<VRNJ\7IS=[INOc61<<CZ@H^=Wd8-g@1dWK.dML1HN-IQdK,P8+C>3W),;6eb
XBI;V2CJQ^DYZPPE@INFc.[Ha8?VI+^^K_#945P-HS8LURN9R&gU=\7N+@568fOL
5#W>_5EMOg/d2g/@<F&Q/3LN3aRVFTQRCT;0K,4ZXG\C:=8,^bc]XAX&M[(=aL4>
g<Ob^>CgHF(HJ#c8P]G2QLY\-bd0RE):C8R<IYbJHIV9g5b#7XaSIST?f6QDZ4M+
IXW-[L9]7M8c@\=fW(E[X+33TV#/7EdB,eId/f0:PAL4P(_6:I77Z_3V&:()I0:E
ZSY-IZ1.^HPgYWb#O;ZDM^\J#\Q;^Y[JM1IVc)<K;6.<^eT95&^O=KgdW^cR-[[5
J@U2If7)[&=XREc&QY]agY<(F82:UOO_TWFLE[EfBF1R(L?5AK]Y+1DYCK#X5#FI
bX[a1cE6^dJ[<\7GdTbY&4#MP9JX2E1-XP5.e2/N-3W72@;T)XHBc[9JD]1f/=1P
5?e01eb8F09&1KN+Y2:@O0Fe;I-PBKMP_JC3W)^69@F<V2[Yd\>S.J-J<dA4MfHC
dFN>a:)D()#-@V->PIY,N09_]Jf??QT,RF?CB_R<V]U6Vef=WcMP?9ePS11=C.13
9_B&Jc:GbdA2;[\+fd\BJ/]1B5VRO\W>Sc4VbZPaB5VZ2S1M86>PQX?a3Yf@[f1B
CM&K\]E8;8DM<6DBTO2ICcBa\-WMU24_O?Y:bD?<F2I+e/\dS_PCF@+_DTED=-2N
GE]OKJ]QZKP6aD2GMg8CER2J=V?+:?XH30NH1e[G)IGI0=0O&4V2JC>S1L0-4J@3
V00-.T2FYI[LBW@-UeO81SRQ4Hg<78-PQZfD&B5C)\^HF/0f^E_c7966#:?fP&;U
d1B;RN<8\GAI#c/E6HcSd_K+/3#G<&V(ZL>WDId:(B()APe35SO75XDdP8N3?4[I
4/PAA7^K.dT?bVf:C:)6]U26-Kf@gU3XIb=Hf#H@?NbSdMYcDIYg()BFTOSX@c0]
A77,_?\N_8O85@06f/0OHT.Nd[6e^H&DRgS,0AW4>7bfX+eGe4BDYB6I-bAF=6RF
YD/+Kb7O#NgRJ[dR\93;CaBe/<\^\32AAfQZ_Z[fcKABDDI-K-G05f.]JN0Pf?0(
dO&]YZYe:U@DU6c0/8MN#>SXD<[BQ>W0]:4F+09?g9-G[?JdW9f\eE2/eeZ<++SV
Xa51>NQI3AJ5c)):Gf]#@8T9:&9M87MML8=(6bf]./fE<_D4P[cT+STcGF?Ia)?A
1eXMKS,_MIF.TX9^0F]MFeEg8HJA<3AIcbU&(FJXfLfX39=7[&e&?)F\A4M=(&PE
Ie.f_3L7c@J]#Z3;NAN?f-eH5_e&@X)3H>//L+MPKV&4XD2aDRO:8980HONG-YDJ
9((>:8.K3DH=8ET4-CY9>LTY/c1.de3e>eP3K8XB6B,X9M(5W=<97H/XF8X+[_NQ
04KK-9JN45]WB[/6:dPQf>aDX<:CCXKWIQUK@L,OAG_,N.fQ(\VK?cIZa\b]=5;T
N1L</Q-_0#.]X:G]d8bfcN-8?0E</fKC0(B)&fU&,,CA5O>L,;Yd]OU4V+)2>KXU
0D?f#@7/Y1KKI28^2^0E]a8&^3EDGVc&f,7W:L(WK+#Yf4afTVL5+HI6(QLG/9A@
6VKQbES;a)MF[>R)YVb(?;@DGL&PXQE:g/P->DBdF2827[:3gE+bLffd5O?QG=N#
@A\/E_&GG:e5DZXb8>^3#:)\0V3TI71agfd1E6C^6X]]gADf.4I;DK<?UeXW[:,L
EU?B<HHcQS2YRf;@LK3L(WXH3g3dQQ[W3ceR52I-;XD7X].a^DH9V<HRIY<D(P[c
CU#M<E<E,KA>S:^&QA9)4G?1F[-B/]Od71K.MKA7HE^MH_RB7Q:E63XE]W49MBYg
0O=e@S3^Q@2+KOU5/e/f?WS^A@3eY<EC7]\I:WL/Pg&3FHA+(-1=EFN[HY&U@fbM
]1a3E4-UE_+1()640@R_CI8<>4.;/5YWaJOTQB7NN>PbO\+f\3/7N)8/_H@7JgKW
01<N#da/2Z\Q.-=;G.M12^&W1R[1XL<RAO3X+1O.JT^(776/<S7_3V_<:G\[4_]8
d)>_NF:@HQFKPV[IBB?3Y&)A_\d0Rbd>XWQN2DHV\/=L?DK-^C0Ua2QG/&77BgU1
N0S_,DB.aNH\XaITe(KeDG@QZ@SFEP:31faK@4egMf)=6<EQ5G>2b^DOWRZ@WO==
bBgd1V)0.TYS0M.3/6^O\6:WLBP^3IEe^M3<[XP/a^LSN/6K&T7,PHEX;S>(I^C:
VD^R(d+8I[HVAZBPd8L<20AAHF:8\9;C]51#?2V.06b:bf:4H,a;YC<Xd>QUZ3@0
E<f>cBAWCGIC[\=;>FISaS#XIceT/?WD72+4>L<CSD5U\CYFU::I5@#5ddBKVTR-
-5DO+T7g?QD2C#&e>3=598b+Q)]?4<B;dN8f(.[NL.N&E3S#8:XJgF293c0L+Bdd
c3ZOb#Ta)+,BWD-\,=R1)AR])@)2GG9:8EG)e=5\VCQ>fVB\(Cg56a3_:+/D378Q
Y9,M?F@\^bUN>G=@Y4XV>&D>DG;NW(2QJ9SP5(?cbG_;PB@6IL(FfQ,:dA]UE_QD
cYX;F(;CP2MP#>,J+&g;KbM_bNNZJFA)/;IK8.R4\1,0aV;C2X9L<&H7W#G,OHX/
TEf1GfE&dH)[Z@c\K@8,&7dK5\JDb5>VLHG6T-H_TfG&Z#G-Z#R;;UFBSAKg]0HP
\)7<]>/74IQ7BQT0&?Jc+/X.c[O\LA^/^.E1]4a>1JGV>F]Qe/\0)OJ;,a/LfX^P
6ED10?a0@-61K4_PO^MVTe[5QGTG/ZNBI=Z+WGX^fDDWEG:C5+_A2c7e:Q2POT>b
LJO>TCYb[dE12VV<FA0,?=KcEMYOO;=KEM+)OO-WW,Z)^>e?a4_b352bF7^1XFQF
,,M0MXOUTd1,X:b-#W:g4,7QY9_ZPb?VE<A6e,C9@-A([4Z<\^CWg[23^<F&AMYH
;9c9^bd[d25-S+[V9JE7IeE0Q,75B1,[cYaG)/5T\gWGBCWKSP1M^>=\G),R;14A
UA;)R1a@9V529>3af8GDGdNBWI6gR5WY>=N0dB^[:O9;1,Be1-+@LMWTLU^gD,3,
7<Rb.dAe</TfVJKaD9@KY&b;+PHD(C>?Td50:3RNZ,#_(c/I+#HYg^AA@EH[D\WZ
(K@#/@^2DD9R.aRI_d^K\H?M,gS=.:V&O+#LEc,.3e]eEe9RG3VY(BK2SVD-U@Z(
a6O+Xc)>ge^bUWIaA?3-KV/T5NRX/W<>T@>NH\2OE<V6>U5fdE:=FE5b^.3[1O_P
/4&-a+-UEEXU\>:2LQMSOUg6)N,&aV64/YbE3W=eZ)GUO&;c:^IT/A7VAE45AF24
C>bDb:RPST_3=bS4c3OR#&J&]YcQ?OCL,aO&@X+2H;cD2R5.I,&@cH]_F4&H\^KP
d=DR##UF64-PIa5X(C]L=>+\JLNTI=0JBRZ\C@NOf7UCC[Y)(b#\DF#+OHD^W;f^
0^,IJ-QNE/?)d:LD;NP&.D&d_#_4+80HEBfYL=^^gAS7CefOP9PVQ72+OBbB^BK<
&2X-.4M7g7Xe42,Q_-A/?4][:N(<cbg610]b-aC-_\#cJ:AP?&<GbccY4&H6YeN:
SdO8GS9_S&H9-OHHKV&TSBH]7&W@FQFd3=;H+PQHQ^IG4#@eg#ZQKRaU@H0SZ:Xc
Ig,=a)[\M+GPUfLC^UI(Q3).c05g\/RPId^UMZXC^gS)LgTcY>.gPWO@I9cUZYS-
P[WXdSeV&KAZTL+E>CAa+e@[DO2+:28T]J;.I+[_B]Y6b&[IP\=]\&Nf1--Ie28]
(N^)dbFYL>(S+e84<?eS)[GDI.N-U_;BZ2afZC:S?\I2PTJ:EF>aIb[K<RXX:1S-
Vc3a1LJM8NbXH#5\@&[U-0BDDSaFKNY#U]Ye^TCA@J,9C[H<b=:>TQ;f<6S.LA-R
:=6fBA3HOA\][C,.-@+M^F1/<@?\AGM,XC6:.@[7.;,1eFTYT@W-&^P,H?g_dE<I
62F4ES\XPf[>A2Q>]bTKO:[gNf,N/KLL30OS6IGB;#/03eDD:df?Yd1?BZMd/A#1
;ZW1>_#FTYV=+YbeZ)#dN8\6f\-P(HSCW.88V0M9P7-\f&G<&(Bg0U5L>:/7eRg&
V,40<ZHAV3\7,.:AMAGeDGe28@>Fd,70(M&4d<T)R]EbP#I=DLA2ZMPS(g07=Sg4
4TH#^2CT[g2H+1+FL.M1Pf9-E3B,\g,N^BUK6NVQ,B\X-9Q[)<9M[<H/?E:#_\F_
;GHK1U+NfaT-Ab=8@.8Z0O=D-MB@_/+1g-KEJW<LG=V1W,[+[4K3JcY@N9RL/?<+
L,#F7bU3[AdEC-3UGG6=ggPfg^?CfNegQ>CePRQ9.6GCUKZJ^_;_eY5VU1B_g#8H
dCYSX\ZOD-N7>#Z,8\b+:YG\cV9Qa\AH6_PPAb#?TgAf)UR+VgbIET?G\V=8D,2e
WW:AOC8@4_&Q+7b?0^eGX0)#J>5>?IN]-)a3:<5).9QQT#Q>:5#.UUg@5S-2UeYe
O/I<V^HS8TZQH[+WG(/_5=ec.<K4GB1d]02J.c5K;[^-UJL47U/d.;gb?e]-HbST
fG3eL0>+T=KU[58g.)CgWaD[]AKHQ;gZEdG\;H4U4@G^:,[:(gcdL5XOLg#\fM6T
NLJ6ZHJFI85aNL8QCP@WT]Z=f0=7c:COSW^Uf<O=?5U6<B8BJSN/9W@;\cG+0P5M
C@08TEBXL;d>Le\6>dEEE^D9B[.>0&P>)^c?#-V@7M8a\-U.4HONe?0RZ794F)F^
\2:=EFNCY?O8>I?;3ZdaF(;OG3?89FHC^[-LS6LSg?@O&7La?\)S(0-,YL3A(+P&
<V(=.Yg;G:.AAb&VOR&J9-:W^>YM:T(Ma=MK7]6#>=7T3f_R3&+IH4/32F_RO:2:
@??U>D2/Gd(THADH30cX@^_=c>=#\-<#P1AY6OQ:AKXRf-YCb#cW@b,@O\T\A\Ie
XfX:V=;]7<<N7/:bDQaD]b[5@7WBOJN5E9:If5aJL0>RZc2b9fDWNb44[(KdTE?J
?OMF@U9Xd,D=dEAb\DN#2_/3gfQbQ6Y8MQP7^:&T3N9:=Z[NP3[\7(H7.XQ<[Ib@
?C:U3BE3J-)EYC.A/^]6IY#9=eb#7J)^fP@T4L&K(ANV54LEcg;BS:IC,Qd5&-3#
:Se-RN0,&1/=[#S\PZX/WQ\EdN7NJ#3B39Vg4AA+A]FN<<g[-O=73.0<gQO_+a2a
c<d26MW#9/cW;#g69QG)#.(=g0.<S4VEEJK(J)eWaJ-\AYaOe,,0I3\ef=4>@PYC
1:8R[&G(3Ee5b5Y=JC&?#eAT8\J#O5/-J=S(9c<2I:PC[)/<Q0MY;C7gN&,)Ba\J
VW5?->@260H0&K@cHO:DNUa./>]<cEU@3IFK,g9WVBM\G?GZU6?f0DJ8=BLa=T/[
,f-01T^W<dCANP[AIc;[eGW>Qf0^2a>_R1FDM#[QX)eJJ;S2EM[UZf(OG2Ca()-c
cd-8JdA<PJ[U2WR42X>O0cHF6&I70Tf^,4(=6/8U-8e>OJT+g#f_.B?0QZa/__3(
ES/cc(g/M^TK?AWV>VL#+B0AP<B97ce2@5KV1Y9E<,P2SX:N-[b.<1X6_E#[a.dd
;1CWDG6D>GdSeLWgIK2a)WG2DHI:+SB]5c]T1KQTRE5LM-N:??A7BB=[0aAA)Oe]
g,]S-NaD0dLbZ:0FPR4U[9&2[?.+)2(=CE9MC/E]RFIeVbD5:?15IZ)E?81\cE_^
WK=&WU8P5b.I2_T1[a1(W#>W/9fb/S@c3NI(+1JaPfYR&?OYf9=9-MG&#>5R9+Tc
P#L8/BF./M)B8F&5PYZf-P1EE,T5B#P&&>?Q7Eg8Pf5;0-L@ENGJRg\+U20>3F]/
aM2K6d-3X.2XJb[=4OQ/N@-a?aXY9cMQDbW]+^cW69Q.H)O&WOVeF@c5Z=HYbD34
JdY+BC&WQ,_X<+6;U;:Bgc;+==;bM)-ZN0(>0&1-+8J4DHG2_f4;-Q^C:LV#Ke=g
4^\O4Lg4KG25<CT^WGIT3Z_.5[__TD=,K:N+aKEM>ZAg_EOFfb0d[E13#>C0XF45
Mc1I.Y[C\5WV]/@B.UYZ0.#(3?3a9=RdT+^N3IQ]bU#PC6SXC\-3M8-cI=IAfR6b
f?CXZ#TaQa;SGY.>A6IFQS&\J5A=52UE?d>(\]8Q>KC^5DdL@E4?=^=ag22Efg_g
1Hc>ZF9KQ;;FbM:L+HLT+I2#RT0EMH5)F+JE@e59:;R?KC)JK\2X+.44fN84E\57
J;[SZV2YM@/Kgbe&;LK<ca>#:>__MN5M.GZ&DH)Z8+Ca1a]I>4f=<+f,]fe/f.fc
>.0FIVE_>gf5fB7.S8)/YH/EMT]^Kcc@<g]CfZG.&>:K&0Q[J>e]adXWHNbRUMA:
1X[d+/4g&X^Re\LM:/@>X6Mf)BU5RY0eA43/Q;[8&6HE;^]<5ZOEf+gId=5@Q()^
B&L\(aG[eTEIg?Q?:__4GQFF\HUgZBWge.bGYIE)A8?)B7D4>S6[0T3ECE:KM>>8
#9aL,H\2.F<d:f/L,eWfPT>L_TP3e;)BD0bSRF3DeX^@_)L/0.^L.+D<I20G8ePb
TT-Z24.eU_HT3g>c39XIeX^(3HLR)ZVJ4#_9.CWU?cS]U&HW[]cEMWU5;0J;;,G+
YUT2K^Y(97VPFVQd@U<^V_c)F3SNd-=(-@KFHIA;bW5TZU;B/bO,/6YK=W>WP<bF
=V2J:LfVRIbMJZ@1fVDgEEO6(Y5-+.[>5X?43MD//4N:IV[@VeJ.BQAd#)?6E-Be
6gd<S:gDU/Ce.S@Y0G=W9+LZOZ?2F;WPFG=D>3.@0@0<4:A?>c]6H/RCJcEZf]JZ
FNK0(J+D@MS/D^4B8@^3PcLXc<f-]3,<]F(OZUK(,/ZM1HF^93+QI1M)KJIU=8L(
cKWPX9QD_<\T+X9Y_?b&aZAA_Z]>][8?^,0G^/Be-Y2O(>(5T3GFQ6?7QXQa7M8V
:G>8bK?NOY.RZL3Y1M4>G_OU5+[?_:;G_DA/;BFLT:@b)ZJ,U/d^3^N>,M.L+ENC
,MPOO-cY<:5VW3^(:b7I95LeYXLD,P)f>F4VMA,/-T\.>Y.>)WE:MG?6IE1@-/YK
-.5Y_gS7#DYbgP@+JB1TgIR&2b9NGUKMgQFCB#O_Ye_gU+W.1L&U\,4^AR<1BI@4
/FVc-=S^;8YJV#66CaK0X#]O4ULW-S>,6XBVUd_6f>O>+./:V@aH^4aY0g+A>PN>
<G4UAV;2;0KgESIKJ4RM?>M<YA.RF2ecIML2;5^OHQQD0e6D9NEEP)PC[,NOO@Jg
,B)[N]VF405M^JdI+^-AUE29(R.@EZ0(7A5gg/CfZ#<8@BPL6=8W.][(<g2cTE[G
0T#5?e=K,7\AME@:YP8F)(:HMYWX9<WGGGIHCNJCE;@A.dR[c(JP3WF6+Ne=4b;7
0bUDNIL[WL9-&fYUNIF5<?YHe[(WG<(,KIIG.Y^_5X>+f7ZNM1Q>RF:(QD?eLK5F
5eHPC?CN=D/>8<RAG^R#;+N363[_LgFJH4,5RN=YI.e:W;BdB9C;6EXNb7c[4P]=
9AZHSFVVEWA/6?27F<<,@>)LF=F?7f&1XU)c29PXS3.<BA-/Z]X8Ca_<dLB9)#NZ
c?8gfQVW[cL8,3:H9XD2HRU,B0.T&dbC)[eb<9SSX^#<c;^3(OKP_)DFgeFTKa?O
MI]K>b;F)]8LTMLYC#AYW9>/C&EWPa>C#[]LL&MgXg]@g@2,P+gQ^(0CMVXFA<+9
P@O2g=88ETe]c4f.<[U16&E8a-+9e,)OW#=1RG2(Y,HBHeJL4WJOC2\6)VF(dEXZ
@E.CY0V3&]^A>b,/4B97__434g-IUPX9&3G9:<eZ/LcLJ^)VPS@TKaJ&&AWOd@?U
bM-dBUC)_Q.AM-(WT\a4UMeSG,H4IKYSF:RT8(c(2:)7&77ZC9#SEZ(YT\\A;L4J
K-T?IF2P]EDeagJ/Nab;\eO4.gL>Pe1JEA?VOV5IZZZ;N2YIQL];^-7JH(^(_:Qb
HY+:DGUVGTWR\H/^P)NLd_[.[OeeRf0<T==EIbQ?(?7O;)?B7e9O7LL;3bK3T[E6
\-VSd-fc#L/_L0JX7^WX);PK:GdHN3eN/Q9:dcd)FEd;X&X:DG1<e8@bbTC8^][V
gMfM5f@Q0:+88,T=-Q2>fC(JHP#bM+QdMSOJ[-G(ASEY:IKb3#.fg2G66H?U:RIa
,cO.T9:0d2C/AH3W5\),=@THFKEB&E#Zd6BS+.JDMSMQKH01Y//ZL[_PJ4(7(NN<
c06)&OQM7/)5.\&cJJP4(4:GAaMPY1=AKO4+(XJ[CUK34e+K8SNX,BNH))FF8Y5;
(0f^0>c6K4G1H]D2\Va4+-@1U.]HVMQ[/[#,+FS9H;?=0Y0:IR>^FM1NVB1,FQcH
eVNTO/<I0,S5SY@&^/@L[F7)IMR-)HWUFf9)66YRN&TVTb\Y7.0M=aA5W&4Ag42?
B[D(bK>=J)=:U:.HC.>SG/f[L\FHgZP[KIX89+;IeEcQ^?(33XWNH1fN[B3D9dO=
AO@g_1]LQg1^4?86R/G3O[TWH]1Z_51.F1T>:g;7[J.O7]Qg7J2DI>P]N+@6cO2g
d@F,ffPP7RNWMWSgEc]=D7VDO\GQBS(YI6]>H9[XPVQT[));dPP16W?UHNMQ/d0\
b3Q8gNKBT-;fA_:_B47b]U(L7Bf45BB=)J7VEY+QM#P@24-WX1Ig7SMR[?/UR]eV
/gF]dC>K5-503]W5<1NX[>H84@_\^C/b-LETNYe5/?J^)b6;A:^;HCZ-d=:Y\eKg
7&T\;X.H@Z9X+),d\:2GM?O,LL9A._A_>JIRfD4M6IB760^^dNa0\C0R[;PNb[F@
+5D+3.c?,0&H/MIBJU?1@(#DCO+03O=<:M^(A^NRA#JKdZ2+\cB5WP,c>3=53O/_
B7b(IB@-<dNHU-EgBX:]PQ6H)=FYZXcR(1/J1WQM?-ff)e_9Zca<R.aJFJ]VQgAe
PF0K5).g4D0JdVcgQ9Pf6#Q\>;[LUT5O7RCDEfMQ7W7JEJ@[?5H#^5,_b3\99MK^
F(_>+T)\:D^3G<VRb1ZcN:][PcKHaKNL=;NJb9[U8I^F8[^XD146>7OVHeb8Z]4^
B6][MBP8KVY).=E<[P3<3BJD4CaAX/<eE8VOb,39:e\8K\[DTa7;#[2^<6IIaAc+
-_X6+2&L98WZI69R9+LK9&g6_]^^#A:167Qc9BI7QFV,Le+XKJABMD]=I6NH<^=;
3N@LYA^OQNNY-LQ4W;HOM#?1?6YV?cgP660^Y]TX_-T#5N3R#+_4@UHg:)O_#P#9
\X\BI>CfdN1f]4KPbZH#0ONNSVZM:D-)O,e9HUSMZbdQQ0W2/_G>YHFGb^2&6_<)
02<KD^T/O&(E?Y.7RFBeW+<8cV[V[badZ\TBd@,@0AYI_M(Y+/D3^+WP-@U7Z_)_
Ub^[H=D2#DeX8PV2([,5?Z=XC;9FeZ1,D28]_cH_g\^1V&/]\U[5Z,dESUU6\+Y0
[5ZA>\(#F_(TB]_>P_eI):e/&?9^dKDM1D59624U#OTZKLVRX^D#?G4FA8I>,I@0
E\4e4(d,UF#++Q8]MN-g57BX@;_X5-)d-0/0+)DK,aMC+S@DTa]93(K?PVcM_/:J
3-C_MF1D+_b/b?Z4&,M#(efe9=YAA:gH4HJ.c-U]HP-9[>5]&R1UfWF<3^<Z-4fZ
R-@,7DQT^:3C?AY,B\8C.;#D4KIcJ08-)2D,@@^BcZ;BG-9@#\,bK#>Od=7VM6[)
OJg=;D&F]H\JS0b)JUBN.RZ]YQ?If7gYU&ABAD=:QGgA=[KQMZ9+bR^0;XVWdOAV
W>MA?_]C-T;P(F;dZcCDN,H\4/NCK,e\aTYMdfPYU_dI7GVgV]Z4#_8VIHc#Xc)8
2Bb]I())J1?Se6WUMcTL7)@b=f<7UFO]PJ=Jga5[Z1&<KIN^]@P>/0W7(8VW2S#E
\<KY55:IE)H8DB3D64.g<3e-R\/MD7d]XT8BaKbg]UKW(IY98GW;&NI>#K&3.J)7
cDDCDRZb3S&P>ePD9?N6[1J(CZb5>N:ML)-:MYME256,6I:V#&)JdabbRb/_2d;R
.a(F9UZWTS;-X3CCU_1_KA9LY2(b,[8#SI<V7(5U#<L2eeOLaPOd:Oe-gK&[N5#]
&9;A_\N#TZbdF2V+&7;3K;)<.FJ=V?C3.0YLc[7<WR50SHU5I4VA4.>X-C.A;agf
-&F5/FA2^[K9S(_BKNbN:4[\SFR91HB;(Y5[\&1P24/58Y<#g^15b?bGEEG7DAQ/
PFX82IR,fE5,e63Z9D.SFgOPN?I.X5@8;NDdVK82f_Q(\QLV\>K]WHS;ZKGRH/2b
P_+R/9E^F\KP^&XE.>W^\RTT:KPSEF.FXB4C5>MC]aV^^G6X4SVa@/Xb;5KcgQ3W
HF(>,_ObM)7bHJ7b_eL&J]#J#;+cg:af/B0e,C.-+;A^e.2?GHH;Mb)RB8D4R5AN
eA/L;02QO4dG:=J#SA<#,4V+F(K.IFT82:@4>:?be&.gNJ[0(OgB>5,SS)HeS&Q@
bP)QdgO<&6U<S..@7^UHe-673ZF]J2gENYJFU+B6TV1;2OTcf<UY_>dM&-SZA3=E
[a\b&b4G/J3(65;9+]QZbPP>JI^GMF<+VW/H.TYSEJI]P&>fe&Zf5[S05B6LZ0YD
HD2E+gAZFMLM8ED?>cRL-.X\+T=KN:X_Mb(e.C/TXJ6O2Ha]8Reb=]0f7:15KEaW
]<bC^RAKM<Rbc,>f3#e6DPBQ[-]>0-_.ZIeA5G;AY8X&YD+-^5T>(6WRf?EK1fDK
S,^+0b(B&E.VS[\cS?BB7d.H^W7LUFaS?QdZRAMED:P4Z2_79CFd2/G>]EK(KO0_
^MKg]C7;Z+@T1+.eUd?@0L7UG^4XgM?e<EW-<448QFe_(FA]=7e3&9AH14\^OgM?
Y0@?_CI\(+/4QMAO\HC#(G<ZEX:1D:gHYK(:W]:CYX+7\JLE+T1=KEUef^-O:-L7
=a0_F^^((]O<-&LaCVSa4HN_G#MNM/ZK)W2\LP@?\dT>Y,O,0>..BYHKd5bZV4cC
1^g=.0R]>FfbZ3+Q_eS^^/XKY,1gW(;W,NX_HL_N,,&P2/352:F0Y)AbZbXAHfP>
bI9#dI>WagDUJb>-N>ed22E4/RVc@39=&J;Zc8d]L>&#&/,QN.,7;5R7FDR0]]4a
[bHU.cVG>5HX1Ff&\2[0-f?_(8NJI\LN4C(V(-/5R#;e+F(G<W[I(]>TLD;#^;ZP
_:68Z]O_fd>3C;IaddRTK1fH>MM<?IJ#)G/I\,c?,\U.)eT]Q(>EWCV=cY7K]Aab
2fW;<.HU<6^,.6Zb2VM,+^aY&+BY8@F[@d-S31f40H=8.2G-?<DM0Q-,0d/AKDe<
?<20[,]a&GA<Z7VgYX4>)bRO2F2&GSa0BFQB:G-QH/RYE.2IOX&2?S?>9.-f(&(E
^Rg7(GF296L#E)S++-QY:=]:^cB&DJ0=;c:917,(3Z85AM06eR[&8)[3//D[fAe0
>D&Z,#)1_?]GA<(5,)X6ZMc[/DKGZ^<)NXCb.OE4/B.+CE;@c:dIb=XT9BSP&.F6
U6c_^JJXaI2X&=8WVBdFaXHRf-Gf=61b]0\SaBPM/;FF6(1d&@:e2O)0_3,MFD.2
XUcTKZ;A/R6/_2&2@_\N@KWc//FObMQ\[]]M1Ce+2+XeC8fBE(U0+XOC?ODT(e&?
)PB:PN)\\B,8@89E9\0X,\O^ZCD&f,7)+_g@c<LfWd4>@3Qb#;,;E01L(_W+CFK/
De(UM)_bYVMG)A;>/K,DOPecCGJ&6SW9_VKdTY>7:7^F?Q:PdG)Yec\K\H#Bdf+N
X>=GWe@9.&/#P9B,512+SU33<7LcQSf@dC9V&EfIKCN_1NeBV#FfN@:FS,)#?Dd9
DK&AX^A7:ac043]?e0::_JF91[UZG)#9fU(-6[2/XFXI3:f#2.@N;1F]MPI=>9Z^
g#WV+-13aEa,LFbN28eOOeF/:5W]<F0/<b3#@C1K@;<PLIPPFWV0H=.:4<9?f)@a
OO^LJMSg;_OAF6Y[J-CH]Md<C\NOOe:8&2Ac2/K0+:/TQ[@b((MK=+.S]1\7<;.]
U]fJ[NF#[POU50g7LB\)N8Q/P)/FGOD5BG)_3@,QL\/c@^9?Z^I)W^G&-2PQME7?
C[E#\9.BXJ-2R3,3(/X9Z;S9(LV8M98U46AN&,@N[M_[>]fZJQ6H1f-A<1ZIQ\ND
JegU]I1-GZaGaZBY58=>J0>NZGbN.4BCFIdB0][3Kd<#4S,5CEEO<+K)7-VTTc._
,LVfdfAHb.VONA;H0-X7OX_&A2#=BH,&?P-];OK6Z;f^#F_.V2N>dNU-?:eeW]<7
3(Yc;=\M7<2dd/JJ1S@/eU]@[@=]&dQ@U708YR1)PU+9^LfX>gQW+0)MLAG8Z/N_
5N#g&C\_7XU0>f;3fHd@51<4&5E_9/_4e9cOGeI8[<fO/,:\.SJZPN1SWY?29@:(
J>&KJHSP-WJ&._4C+T]6eRd-0?EfG,d1:SX09X79;TcTX1,TX&+c+0YWGB[N<2gH
?g#-W8A70:fA44Q^K]<ITed,=98c,N99YN;:-12BULOOZY,50_[)[NFg;?T.d1^d
ZgK;EQI\gDcQ2CF(dUP0O-(Ed#aQaO4;806#2DM:VU?E4:T/C1:ZGY>D8,&+a.E,
d,=C-BOHUAF-CA#PV:YH<;NY^N/HQbc_@W\O)KX5Xg][7>>a80D7PP9=2Le6=eMS
0^?Q<JH5,>g<W7]4SVD+d;O8KdbT,^aOLSP=aD4&@B_9;d^<6SOHKVE_<gU=G07G
CUAf]<21&MOUK8<DB9eK07O2Sf^._-Q[)8GEO#Pg;b7MR;3c1c8VMAOEGDKa==3>
Gg9@TMM/RZLHg(9.__R/#=EeSGTg5C:5R_.]_A?dTJXPf9D]OC-T8]aH,=)I]N>K
]O^dO+)32[79<d\U)QFFeb,.g#g#6Af0VV4^^\6A590Y83[X813CVT33.[cSQPGN
5a4=<bZfG>[20?/+_]W)9751>B9c,]MP_WAdc0<G_HKOYMCUAKXgWM2Hag(@fUa>
9J:--/?LD(A?VN7Z.VYJ4&/D\V6aWQZGa,DB,JCD(D?6U)g9.[ATecFRc_[;gcZY
W=?,NPSMEP8MdS.8]b(4LL-.?Hd#03QQ[)/@8fL-GDaa1,BE&0/\X&fL5]3c6GL/
SYB3DU\dYO7JdF;=cPEce)I0ZD@Z.Ogf?MQ/X9dgSE8F&TTX7T/&LCB#H4g6:c8@
,5B6/g.a4f^L^K7^@KV<A>R5E8dQ/7U-dIBLK_^4K#/>ffdN(+2A9f3:=Ce9eB]/
abXSXU;BF.0=Q?[gB5,g&:G;UU[@?32O;SWSX_&W(0T415Xa0#W_CR_+L<59>g^=
;@UR;AGIPUT8L?]5OH8,/:][)9E(SHbC+N^7DG4G(WEX.AE:QB+(WE6^BB83TJIZ
e:[<a[c0DWL?CZ>[-:SDS[GO5H;8]eeMH?U_g,eGU^E,<^]XCNZ73Sg:;MHa;aa?
K:;&2\@+UU0,<07-MUNB_+2<Z4bgQG<-TgQ:-,(]\P^98?)5G<JIBg4Z-W,M,_V_
[SE5[HgIXgR46IRTO,]Z:W+WLNf?V)H@J\<[M/A(fS.>?VP#/a5)DPIIW(E6M61d
f)Q_?=02PFKND_Ka-DN=?0_H(M;5c9\MSFJ5Ia<3A[X1KVOJ^]1Z,.5dN^^1[@@9
&N8aXOF3_63Sf>OV[CP.30(0,?5@)\beW.6=:1>cNAW]b_N4;:9Y2V>Od^,-Rg?N
FUJR:cXe<--XfQO8_3HB(;T#[:2;+1[L;gcY<A7F]Ke;85T&XeS@?cFANe@Ua715
WY]Ca#.2Tf2-0P#1F<BWg@_X7DfUH+EE@Q^+_XH^6D@#g;6A-d?]1Z0(;/OT+\G6
&8bWLV6bLNg-U4?=7,A\;GY:H4caS6c[&^bY1M1c[S-6-2aR3&G5J3JZ\9OYK^4b
<Y,:8_K7Q0b(Q-^Z28S3:?]YVKTE5,e>TED9E;8gJH_K-:\5>g6-]L3dR:d[#^>[
dWF77_RW-/AI<<OA4AS3=e=IF1:g].e[ZT(;W_(S0A..Qd1a(PA)H:(WgfBbV>eZ
AK7,&40L79?J)(>U1F?5EVYBa=V<2)?d5PV[I:135Yg_Yd^U)^>3e&ae.=44FV.M
R+JJ-SJG-IJ[-1E4RXDYYG9R_T+<IfZ-7B<EC)30U_E^Y(B.b>dEf[Q,3D60=>U:
Y/e@YMA<]6VPHXc1&:B4^0EBA@R]NC#J/CX(H^O#]28].cAN_HVV(eGG?PE3T\BD
7adK^SF1\S?#0G0CAM)7:cIf_Pf:\1LXP./KbC,DeU?NJPK)c#;B\cSVQKBSd+@G
JZEFgAPH6RW^cGdb8LYM22Y-C-TVU)JcRWX&W^M[B77_9g@J=LO5b>=a,eQ=H@Wa
AOKg8d^PA@H/cEaHOES6f7,T+DJc:Q>@3K..K<g/5;.G0_f.VP23-Qd[bE;Hf5\[
W;NMaB8]-@g.-BBNW:62PU.PbWB4I,_730SF_?A.87S4V1Q^QAHb>(9fa3PX3A48
M8JA0I_9)^L>>L^Q8Q,EaTZa&-;5J#&#:dA&(APNZ5EcIK[ZcU4^\cO^-OQU_E7A
RECSTT#E[8FaH._J2^2^JPA:.;_(P>e3L2L@T:dQ/IYV1>#E;8??RIBGMFS0Gb(R
e2-+O&.2&dX=_4HU]CY\^RGUFRR(ZEH6A(bg[W1XfcYCcPH=,8:(-5W2g=gc+=N+
D.T-@PL5,42#CE/dSI\/b\.]7?/fQ#Zb86[B^B(_;M7PR-2XUY&3.BY6VZaFeZEK
RPb=HC^f0-#J8HL<<RGf+Fe+T_a1#C\F3N=/7<JQ(;T.[g47QVX<H73_f4WC[-V)
#gGH-4aZ\Lf)TFaP4?9#Z[XRXKBKAVb?O>C=9;&WKeM8@A7:Z#)f(5#c3E@M?&CR
L>36/8LPe8_\V_4VO=?\/bS\6/ZS7)]G,MQO0Z/G<H;P900bgX,J.4(a;7GJK>CR
^TOge5ENA)6A0[9+;:c/Mf&7O-)JX-X?d,YV2,)SdPBCMO7=8Q.d#3\7P+#?-cO=
b;aff))W/Td1:2VgT2/H6.gQBM];\Bg.)[5UV4a&fHJ[-E6?H1_2J[\4U#G08\A6
WfaSaD]Af[>?MPMF,-RPA:-23D,8=b1L@0/d5>@I9@e1)LZ9@7#78^BaAT@[)IR<
>M;b&EIc;Dc=3dB6Ya1+S&a5FR/eF.SXaKa#Z21UW#1H7QJRATW(e9\8/WB_P.0F
HgL@J.@7@d_Q\<))XW7P#49/JGQWF@9=bUV0<NWKAUUHW\.Hdf3E__2,fK<I_H/1
HOY)&:..e5Y1C4L+W7-+T@;:9UgAP+F/F(PH5>f:_>#]Jcc4Z(N96.J<.]3gFC5.
Oa\XTMG&F[7YG0YbC[]+Q6,RXFZ#VWeT)G#=/M3A^4@eMEY+OGFVgJ[S4(69cDRA
?M/.C+U--bK([G?(Tf=IES7:.aSe.?X2=8f2_W_W^IA^gfGG9U75614B.+)I(CV@
/&(gCd7XL=D^1B-T5:##Z85Lf0F;QA?:OacYC^@.)27<e1CH:8FX#AEbKJG3-=R+
LFcQ.HBf+NE.V&2Ua-EW2\-8]ITMg:_ec#?&YcG5U_/(IZ0>,CMCUTMLQ+HLCHQ>
D54>g?S^eKI^CB].L_bg146K3:dGMO?1dO8P6SY^b_,DHQ8)^dA411F].4>d:[bf
-X=0_15bCBBGC<S/TO_:>88^>&GWgC7YGa)CYa&KT+TCA7V13PDRB#(UJ2?5MX?U
D8LSc??3>>S:[LJ>#U:;(_RX+6DeY_&]@-&TA/S^_@R=G]ZY[HUa4#YG/]a/=:b(
>@c\+Ig5[>#U+T&^P9bL;;6JB6/7Z\;QO-SMC.W5O(CDWV2T:7+E<g,J5WP@5EL_
>VV4?W+@_S/S[a\8E>E<V(;>6E-./H(=-4)_g,\-SP<DDE0QS</KU&MNIM7;3K<#
07g](X(#MTg+.Re)O2egILWX-4DXPE6H67&D<UaG0VJ2-?B:Y;-),57?\_DG(A_L
,4)&eF8>IN0#B/XEQMLJ)YPQJd-W3WH#MJcRJOSQ@L+g+BX<e-W];;)9H&)b6A)C
ZQ/>E::2_/g5c-?S1Q;W[gJ(=[Qc=#[E]GJ7@-4PU(:U-+M\)5KCVA2cQGG[Z6Q>
=?;PT;(d](Q_76+B-[V:<VKQfQb9U:XEGPZJY>E3B-8cA40,H,A:9\OT+6D9[8Ke
J>,(X+R/G/)<P@5g6ZSd+.JbLB/-f2-+XfJJcfI3OKB62/O\S3)VBQ#()XZ0D:UE
^c[9:W-c3PNVZW6Kc7&g^N&IO8BA/Deb(;DbULL-P/]@U+\?LWQ,MB\@MG4T(##L
eV2Yd0AbFSdf.(;B&8N4U2RXd0>FA,O]FNe\_GE@7=?B-IcS&QD1PXTIA#QZI=f>
&)R_Y6+W-<QY+A/&2+H2:(W=/P1dZB>MMVDbP(+,=&P4O5JaeOLBg.5;DAa2MENQ
H7K#A5)P32DUYV>eZbWBWX@C8,aJKI7FEU)H0Eg?<[]:f;5FE1UYb323J\gW&HT+
FMTO>_Gced6HD>1J;<D2/6\:@/N^aNI4e?TN9dMVHf)6<N>)C.+E3/d2O?28GW=(
JQE^--PR<\e74:S_McGC]f3,f^(BOC6>6eLM?&Vb2acUHX(4_<I.4_Q\7ZV/GcR2
<fA_2b401AIg4IO?W,+H?)SM431].3++]IFc]8Kg4Lb(11Q,ADN^M(\,Ze47a8N&
d0Q^2?b5Z,F,4W02),J3X5R/87,VM<7_7QPBLD/bV-+U[LW0KSOBR]^6D;>cJ94T
ET3f[_+HeMbAcBM4Q)U_1IZ]X@[^6cTQbX.Z\9#[I./:^C2E@H?X(d&:-e6<6+;Z
:YG#JKBV#9dW4?fE>?5P:PgD1(.)LG;aQ9HN,0^>-X==:ZGU;9MN9_0.GS?DcPR+
[5B_X+U?,-4]Ag5<PfQO(FGW(;U;7FHe:D:;)+Y;SAO4,GJKcS2_2,KQ^6K8F19.
fYI:PM9H2[.MbWeOXJ#PH&<04MBNBA>-E]3(SWc1YR?>_1@ED=RW;DHU^0[39@e#
M99gc,Zd:IQZ2cA-WR(NHT5V+4-H=F0YU4Z3faXcFT4#[MM6XWBANYDc2R(X1)-/
N&8YGSa:;0R#I42(JP_ABI4I1;<d5ICFcIDaL[aKJ?Ig2,3XDJ#>VNS#4&]P?:EX
7b<#JQFJXaK+M(QWFZa\)aWK_HM?#[UHId#b5TM:[AJSR#a?3).NKV6@dF2I#O)8
/e_1/:10Ug]J+&.;Q.F6MT9@__+@X<dYfY/@[.I891WB(]>D1BHfF/+Pd_W[c:JN
dgJVPP7#7BM7W1VVQ,CKP18(^H+W.@?5X?O_/?4+4N68KEO#K(X-W@FQQHN^?_:#
)9FY-bEUPQ278568OV&R\IEF&)b_CGTR>4IYV[P2[bUDR^U-B?2)?.=07g]RLLPE
9D9GF.YGUW1cIJ>Z+e>KEdI4#1aUOgQO,Q7.UF-P6X&aJQ=8J54E[7),D6YQYQ=J
<@;_CE5G0PZT1dYdA<R^AOZ6HPf=U<5#EH>-BDX^<cKEc]\=[U4@[cZ1WQ/B]2eW
ZF@Cc.Y31KZ=66HcI\NgK\+OHdZGVa\aJ^QHf9AbE^E-7.b33@S)7R1W-]f1E\CY
F3IJQ.b2?aDSgX1[#?R@U]N?55\97U#^JR7EcC6O:,XGLTXc>UJ+d@N4=7NH=(df
C[b>O87UZA/G^Y181O<[a65XfXA/^<P)6C^<B0aPeb@FLRG?XXK;c[2C+V,b&\eF
9,a?5SQLWIe-^c,NQL?]\1&e>?.)eS)Q,dS?Q@^g/g7@SWO1b&D7Q@7_a:M-U&3T
=Fe.B[b.M25Z0Ea^M(1VPCH0P4[98/R2a^gB)U0bfJ6ZdDG:2>O9,1Q-5MUD+g(N
[Bf8UP_d-SS4/L(48GCGLB@R8SJB6W:(MURG91=_X&:QGUGI?Le[>8SWW1,ge49C
VM7P/X,A(Yg-,;<b6E=0A]803d5)#;U(.2I9@[6f;gOJ/VA)8X[Ce7CJ^&R9YTcS
EH5d3M+5dgR-7=M#dgP16LUC.P(K^GN^PV?,M@+A#9Y/G03T_R]=];.-8KJ-\#R<
b9GK,HK8HKHH@2Fa<QHcaN>ML)V6f@FF7Ob0R_LV.\\N-(B6a0\6TZcD&._ENKRJ
]_Q9[O91QdfgNIV#LH/T7C:(MHDXC9>9b]1VRS,A.U&W#YH6(LbD-L@Z=FJHNBUe
b=G-8WG<PBXL>b64K+DXH>AL8Q)ZW;@K#>gg6dX-bd9<DW72]G00fVIEf&X0J-0,
_[WL?F\LTLId=ZL&(dCKL?K&Z8J?SF9RaA8MV)_T26aNNGOQAES,b8:-Q,N?aTdP
XR;9YfS;C\eD(C0+:G^O?;GEAK\FD6Ha)FXYW)]=KT=17QDR;NK6+2CZ#P-b=YAf
Ua;9E_WPS))>8c3HIg9\d@0V(2W_-2UN[.>T9,.0U.^O7C,Xg8^F11]0Q(Y9>b_<
((83&S@c+:I]f+,SN-T\gT\cM[NU/J>d5V,?V)3gLPCC0SO8N2aR=c\Z4UE<L/ZL
?LFW4^;]e1_OIB?)\1?NY).>@FK7.25a9-UX7gU.=>]G\TBb,M[0)0a>UfNg)3W/
\+;Ld6ZCURYZ+H;^09UfbKK3R(#UNKcRO<(I?,FFOeF_@)OB_d;UY+42@]P-J1?M
U5GE^I]P^b)U0JQP.g71>99Hca+BMCa(R+Oe(6T&HUF+WaXL]W@6XUOW#QfbQ4MW
B854RUG;,Ca&#EVIg(fKEJ.P,8UPdC82CbEb+.(9^]PQgb@B,3RAJV02J-eAWYg<
3PHDO\\Db_gWV22\R@_):+@-2KScNPP75f>&VI5f^Q6dVDbJHBNI,QZD.Gc2R]-/
_bJRNEEG9L=Y4:DddW&&U/U<L:CN62N#2d7-MTJ[cbXAHObVGZ]f9Kd_cJD=b.M(
M/6_V[AW;K^5M0QMf5.=.8)3dW09M=RcIe?CLJR_fY?WdELLH7BJ@LI>]_-d.:NY
C@R2@G#VgUP)Y?TN?9Fa#F=0^H3@@bbZ3W3,U9;-]KT(_E@X,7SSVV=/S3RIe,L4
UO7QZ\>AD25P2=aX@)W;-G/ZaV<OO3-CGC@;=^[SM5W-)?Jf0d98+FQ)V,HVKPQ9
#XObRDGRCUHC(GR7IUfKQAgU=\O953:J357JBDR:?D/X#X>dCE)2P2f[fDJe#F6&
1;_T&9A0-d_5D=_e;ZCT+)L\J7?=g#YaH5I<T.TT]f>0gc\\J+@^EX=8Za:KLN<-
OcQ_I2I;e:R.>a@d+HNV@TYXf;DM=cO92ef@&N>T2(>EI)F\5W<A^AeOF<ZG1fc5
Z6<.dX7YDF[+W3>]NUe4:9+R]@IJ<_(F94CX,:B8?OC0D-F_W9X7J(VcFA^_UL2>
0XaN5VJCA3a)>eYX-B[.09P(.3S9S#-C]\Ef+A[,aR6(,c>e&FHY8[R]&+UVGXI3
R+4cE?O764Pa88)F8a1WZ#eZb0FPTQTAY+bKcAaeEX[B=\Y:,[Y<>bHd&&FDS2),
d=a3e?R@/#6Z,CE6H,\5#77@/UVVBMEX(KRWKLD_-/1452-6,GJa\81a80;9#,1.
aaXgMNJ#9B>CEH3fE-H:DEc<P4<T-DSRGQ@>+AB/,FdG[(MER&SYVY)/F^:M9CDO
&:GOQYRgGP?BMA&CN0NI4+0XN<0=_1N@CW1cL\OF@&g@W(O^Q5.^,5[+0+FLX/(d
B.EaRNC)&,BX)E6UF+/O&dTY8cCMa2P1>(O#\/>WZ:_23fZ&_9cCR>?(=?P^F_:J
VS,S5Y=,_R&IT[EE]QX7gG9HM<ZLIR\S#.+><:VBACA(MPF\T]b6CV7BdR=#eMP=
8FYPM]+:E3M[<=U<Y5[I\@)A\gJFVU#dD/;YC6HGY6,MRfA_HaXKa+-SS@A:V##R
+#E/[K;K3DI+PPdGQ\D-0#dQ4?Cf6(.#IgM;Qb4?S0K=3J#O[R)4cfAg<fW(=Q;C
;,NBS;bbGBbd\-#ea(?Zga3+Z@ULE-ZAW@&65V[Na>3Af-I/Y?d&XQ:)]\_f71T>
0O2V6JgN<KF@XX=9EdZaB(B\]=_B8@&H]1YWA>F)Wa3UHMD-AgVeS2a-X.3G>G(c
L8:29adaf\G<)TR&0H9\#M,31^F\ZTT&bJ>EHMX<(4&Oe8E(ZcHM^:-=Fe,PgO:N
PJOHASA;]-5e@D+A..7IAO@TXEdKbXO^c+U/2S3\IeAU9M&F.9PgPRCPW2E:D/S>
UB2ab],<X-Kc,+^6aCM[bWX>2@-Sg\&>R[g):-a89^+[V:)Mg1IWRKU5Nc?fRN-,
fI/DaXSce(E?+HHW,9a^=JSJ=<-X_gU:<Y?]^+12O9bdPGPJd\[SHE\@:Z5##@\5
>.N/NA12-GHe[DT=?WW]]aSJ5$
`endprotected
endmodule


