// TA demo Pattern~~~~~~~~~~




//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Siamese Neural Network
//   Author     		: Jia-Yu Lee (maggie8905121@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      50.0
`define SEED_NUMBER     28825252

`ifdef RTL
	`define PATTERN_NUMBER 8000
`endif
`ifdef GATE
	`define PATTERN_NUMBER 1000
`endif

module PATTERN(
    //Output Port
    clk,
    rst_n,
    in_valid,
    Img,
    Kernel,
	Weight,
    Opt,
    //Input Port
    out_valid,
    out
    );


`protected
L1-@.E8X)&b3FYe\-fG;WMU[W?]S9T[2Lg&+G==G&5/XFDIc6=_U6)>:CT;X1g#F
(:E:aD56BMX5PaCCCa4GI:GLSYA(dgJTIa4P<[,PY@0>-b)=9N\[a5YC)Y7cW^-[
eDN/-Sbf?#8b>SCPFLTGL]:(Ae:2X.;)U_fd[d<@dfH>XVFfBR-3NI3Y6(_Q&,dg
OZ5>.GN#L_4K9JI8F?EeTWRI#:CR9POeS9QO9cSJB5]QL;D:@25TNRFTA-d5NDbK
FHD/bWWJ;.IFVSgdJV:G(^P5\b]O0HVWDgQOT7Q5IA/5ID;R>_<d>9FTK$
`endprotected
output          clk, rst_n, in_valid;
output  [31:0]  Img;
output  [31:0]  Kernel;
output  [31:0]  Weight;
output  [ 1:0]  Opt;
input           out_valid;
input   [31:0]  out;


`protected
+Ra(4_\,-5/.\Q6D=1C4:DI]0P6CMd.XZ5Y+,fWcWC+C@=+J9,VK&)62?<>MHGY/
E:5Y&C0IKZ?/gdO=SC5\aI=415#.>XJ7L_2e6\7K\IMA&GS_Qb<EgJM4V+c2=4\V
U6/LL@Md\/(A-IT<LgTab+e5b,/[9,^=Q>\I(?bX+.+QN75@;1/7c.9];WI[#1X(
a/OQ@NH]4ANIQVe)BD:NDb#H;b1e4TN[<^#P>YOQMPCL6c#7C12X5HPD:2-Z,]^.
5Qf#Q,0;e-0ZDbF>0A#HaBIS77K>QF;NNC.bA)e0:^bE8_@M[F+>c-X&Z6A6Qe_/
0=C?5IG<6FgD+TaHE5e[6\K2X?Mf:1)[Dbb<_JLc:?\+.,4C_+7JGQ6(d;Sa4Mf>
S//9N#,5LaTY^J5f7>-g[Q&GUCbe/2Z>._e(BEGE+6XJC@3TfAT;eE5U[feHYb08
[6O3C\&N(dJ]J-b7ES8D?A^Sc>J3UMNDU8FU#]:^&2<Df8-ad5(E>Q9a_)9Zc@=8
V6[#Q#LW(T2<eQUR-DWP&M@BdcX3R)PDNXeIJ^,1<cG5B;PTFc#LYYUI.HD1,MJ>
(VD2dX27:UK[+>BbREZ<HD7V^G/gJ0_C:)V>-5g/7?5^DHg<f@LdQNb:/K)Z&LJA
,G_8fB(Z<T<g/ZUeT-5DfF?]X;8HX93bBf^]-P)^@D-fEAbX)&)[?2TGF^DXB2#]
K\:+=-6XCUXDVCe>:C-a4M)&bKYU^/W.6L-5948;\a\Y,[=_YY1cL^W3=><cA][[
a&;/UFYY;8WI?ULM;AeaH.Ef:):6Z^VegdN31)\,8XFMR31fa[FOB&.3B]c#U015
aI^ISNB55;KQcO.<:E+bMZ0O74EM,[4L:]af?U^>U<K:_4U-T36Q,4<\HH(86TQ@
][W_T49RK[\8e-.YSHWW@V]F2M+7>b&=FgRc#^a^<=\EM3VI3Q+=_S:,(_\K-gS?
U\TU=GXX0d3[TZEE4dZB+OBURe+.OH6#4FHJ8(XW-DNc.K#K0A5J>26-W(@2QT\S
<JB?eM49WB-=_UbDT@b.#=XQ1g[><Y.Vd#LMPG=GMW6N=]_3;Z>bU,/?EGgSHE8J
9VSDIL5#GQRZg<L[-,OMEX/[?fEH_PdB4VQfGIDY#C_0/BB&L5=6GEf.f)F>cR9K
@DfgeC9T2&10<dc+<7-Z)5g@6:5]^MZ:[EAJ@0XB8>2@T,R_,:GXRK[DQ]fafVM_
8CaX)?YW//:7:N5FbYdfRQ0L?BTB:Z@DAAR9?<F23K<;(#b^GeNM>d2R+I;[.^ES
=[3GVG4)fA:_9a)=ANWKL^c[8eAG)/(I(OZ(70:CN2L[3K\8LYae;:7^/A7#CONg
ZLT#(a#)S5ZCZ<?5:TFEYE2-,3\/.@<]<3?8^O;(_M0R5fKHGgJ]^IA8//-^d+AZ
FX1]d2bGSZ^3.KKEg8aS1D>J[FZ4TI3G)95<5<:GRR0H/B0XdHSO>XV>OQZ(+N<6
)6+egg\_6PMJ)Y,]F/HEG(5(;C,WHZ(_XU\?V4Xb0Hg[VgNW135=O8RW?M40FPYU
f7.W&eWD5GXE&D:1QGSA-;5C=W\YNd-UgYQ4?X.A4BKL@8[/+g2?XKDda?UC75:P
WI9H:(2R#4A0]RDL.BITg4-0a[b_OD@6.f0IBC3M8aKN##A@P6c@DZBXE1:Ha>&T
4<PcIFU;&V\D<KM#<<VE]0>37)&1+X_6))FV3#W9eV42,GR/Y];Ma>Z3J-14NNDT
9A>Y8+42<:QIIQfLV@AJX4:7#97+]U>/\beOQI)CLe^&\+fJIAd1/+W7gN)C/BM1
H6,D-bKK.>J.XJ5O&9bdeH0NUbW\QVSa&bIYecGFE]JX172HTA.^QGWZ^4PVFbZE
GT^9d/L9RX^5)YJg/>:\HL.X/L+D81:.c8SDI)<b^=Q[6W-?GSIa_LQBE]]Hf]0.
;Kg&Y-^2<X1X,+F6?WKEOL&OZS9,/\4-/;>>S46d#:C=PIQ4Id_;UQbe\RCN/,NJ
<=7:gE8=aP00O^#C.(7EeJ/]7c1aSQ,]9B35EgGM0g4:JYO@ENQM&54U)WS/GgZd
f&_1d<aDWBeaAKQ<_KWOKT>94X.1[N\1&>[?<e^ODgM^=:fE8<dRXJRHPf/b:+V/
aD,dDZQbfP21.H2=PTF&3;.5:\gg8QPJ#5S;U+V@HUHEKDL#O5D5LEW&237gE2E8
R?#_<=^D]]1LM;P:fXM77H05;4B))VM]@EL:N^<_5/7:_+/0I3=.6Z1E+W88LA9Q
HX+AH62I;@@1aNeN=PR3)_38[M#J:4FF78)+XYEVgd#X^<(bW;FQXYfR0LSA_PQ6
>A.bLH;db9ME0FTVJE>8e)Z_3+TD>.7dVY=@MU80MZ\,TJ3U#HU@dS88+YT7DOGY
JUCC[1(FUU52@7eB]<\,\)YGPR2NSHdD;R;RbE1(:gRKW]?;Y+3b42YMJ4+.b6;E
[V5+P6Ga3+5P(+I@bfG?,cDc13e-aDW0L46L62UF(B,;7[^,ZGa(N^==ScQ_.b9.
,dB(.NV@CIbJP8R?_\PC<(IBUNI.P4FcV?3ZZ=<65ENDGORTTH/b->?L0fdFAW@0
DB#&WeI2b.#,5fbMTGKKXFRc\+TLW(c>)WDg;gC5;]^I\0[>N=A7#1@4MV0GE6fI
O]ZBH0UC4M^5<^H?QJeE1V_4CW@Q&97RYJLB;LX_eF-Z7K_8>Z_#I;NTC&MW,J1_
VeNHAHY)AQPW]\e<Y+aN,SfL3LV-<b\d?gKDd)#<//;G0&@R41.^?SS_IORQ6BDZ
97E7aMPW2c5=5dIZ7[MNN0O7+V)/3PF7@#8,4F1eC,;SU&58Dbda73fS7XYgEFKF
E_22V<6[)P3>4E\;&g>]G-H&Ud2Y]DVO]<(U2Vac5VN.Rb.M-,af;&FS>_(<Vca/
-=-cMC+ZIC,(PLQ0d54G/VF1<&Q<#4V?L;W.CVA<3R-9T)R1]de3_af)]=AYCP]A
>5)4+Ye1<DCIa_ZPV-@TOM5>gdG]BZ9&R17:HC-<c,JecU^B5BOSQMVNQYf0YV_d
H;(@-T]>(](bY3,F4M.-=KdTeWAU.9cF2G;A;KBPebB&G\V^W6:#S[68R,2->c5R
W7b^BS0A[Ac[XK9/>_eYZ6Y.S4Q+cR#V=bH_60LC7gP-&]^ML#J#?[cKG?bX)]Q2
[?QKD\C>&QF6)8N5/NccIBO;]R-/HIMfBKHeT>:)BM@8CP]-S,C&GU7^R1OX)\Xb
46:XbRZ=@J2BH2CEdXPPNH;^>SOWKX65Hc(@O+^(MOWBS5[Zg&)TXe#0#Q-N\(D5
DJEV3:^Xg8S9cZ)Ob(4Kg@)g,aW@@(MJK+@O89&3?#9.=+0d,^;XC2AX:.5LL](^
-ZKdOK7JL##dDC&165\6SY;eUTMg0)/&6Aa<M\b7>:6OH&V2ZF;f<BP0eaY9gY.4
DTE40G3=ECR8TTG@KW9dKST#ND@PRJ_-1J-8,d&4FadOG06TB<3KHT7<9-Qf&SZZ
KcAD/:-TV(c>,7P<>>;LLfa]6[5JC./^80V2L2_KLe7SAWc+BbB+g=2/_dY1U20L
76[(2M>aI#FO>I-c;Z=P&,K5Q[W>Md(TN2]/Sb@XbI<H5LRN5.>&bW,JR88^8-9:
3Q(X:>)MY^FT5M.eVAWb+ZCN9CC,>QIRT\KAX]NSb2:5HE(QXU9?R\gg[E>RB4+)
7>QCU4IA>-?4YFaCeR)/&J2.VK_I/ba9Ead]?a4?2H53bUb<RMD@RJ;EY+3[-QV4
Z7APf>R7<gH25ILS^:G\QW<I\\MGdXQdUac.K#^f0R,O3[NcN:IN?>JVQ?-55>gW
TZT8Ud0AVOb^^/^/.;QNHH8W:IbgbK^fJXJ=1A[<.:e5>)Z_R@0[G+&EU),YQeT-
6f#c#VUJTW?3]JKXX;9D?T\?5#1Z1Yf8],2)3Y^WFVU=cFA.SF7C:4IK,FBU1_U#
4AV=FGJ)M9Z\eCcI?ceF[,aB4)KB2H(a+1DAMeIC^&aD=):b-C88<]EL92+^;Kg0
GeIK^(L;N/4gc5&SGQf<]36d\[DLE6O,0GB]ad(Wa(+f8ISOEQM<bAe8D6fgd?gA
Z=D=8+E.(g9WA=+M),7[/TS,T/I(@1A90EKZc,A+.J@0>.?d[&;3<\g)WVOWW&5U
PL.XMQb@HdB:B;^K@-@VLYGPUDcE#LLNU=cH(.U9gFFD>)2Ne#NG>7=Q+L(C?Y5P
UW5)d5H)VEW_9&6Fe=?bG>2=.fg[FG4?3d>9U)3[<.)a9?G(eOd\D1bH7LP2BeLL
Kg#A5AJDP,+PLYT:[Lcg4=6b57YCFKZX-V.9L:3:BKeV_\=^>@?4(9@Ef[)6-.TV
L>e3KF]1Z@=#A\CC^7&74,]6=dXP<3Kg#E3WSOQSE@K[C(Wc;@eJ.9A#L&:&E+#J
5Af_-]Q@I69#_SN4OdW7L<#K5E@H+NcQO1,eVOV\gZVUV]2c(O:6?1C:]8KC(]dW
0\-C+&D29+\5Q=HgCb+fg4EM6UfL4EFH.OJ<SdcA<FN_E5L.5QfCd3RHRLHgK,d^
-@54CZ]dT>3/8E^=G.#6-375BMW8S^?+FI[K<?D:O37H\WG(M6Qd>ZYKPFVMIE2D
RY9d&6FX@U;ZM3OJRbB#1HX.gJRP6RH)A[Z07UcW.\5W?15e=(IGUdC+?]6X-79)
,=9;JQQf?F0\PPS6_O_D6Z^FMa6YQ?cGUUCQ;X3PP,fdc.PT[Z#[]:6\PeHN.NIM
5TfYS1-;Z];/@(QPe^.1OfOfYT.K&CT0\[&aHV<54_DbU3D-WUJe^SbcAWd+@TEZ
_Q.=5ZIgR\RcGYK@_YZd\?DMTJML^bZ5L<NW7,(G-V(:-#Ub_LeIKR[WRIVVg43(
;4CXA^9?2QETNER[T5YB>/2\>IM^>Ic.&<<KF)67B>^+eBfP[D(NJc-#bB.d_Y)6
_H#8FGgc\[>Gff)KD?8^XKV_\_eK?;Hc,=81;HH^@BSC<(7;40E&P:;?+c3#+P6B
=Cg1MV<9^O8T1]T)2P90XLPUZcO4;d8#P&A)-8(Z#3YDN@@AT68TP07e=>PBYE4a
?d564YLW&0W^81)2VG57[PAgEeg@V^,gCPZ=bd0]0_6#BN=eeBb&RQMFH=50?WeH
d0(75O(RT3Y[M;)I(NEW=TA^G@]7a]^9L:fb8EIQNTP1M7[#Y)ZD;V&9(5ES:JbD
_[Xc>)9]Sb+\I<c&6<Y(Y?e8cVF9,PK](gMZR/])_DXc/2c:U-N7MBDGF3Ag>@VR
B.X+2f2DcE,5^F0YQZDX)<)[EdA]TZYIZK,SGaYKWgg0VM2R]RLQJRA+KY[FEfJC
>GV/-.Ug1\&X(c-53N>MD(SI3aO0A(.V7W1:TdK-:=I5NP23dDCTYO]:Pg7202eA
TRXHI_eY?g+9dTG8E8<:B[RT7?JXPB9NT(Gc3:.eYZ.)a[M9CUBc_\3R0J.I#d25
,F34OD8MRcZ^@K:?5?.f\+WHEF6=ZUT]L0VHf\?)MJ[\Z;HBNVNL)+-MG>B25<CC
4WEO_CH9O-9E^VH_?\<4[;eW=FLH_]@X6d:dNKMd,7U&X[TBbED8?]PGFFS\C#c2
)C#LYeR^AXfXVO?Y)N&7b?YHgg<e7I:ECE;<H>FaNPZ,Y2=5@-AOCA2gM+B2(c,;
;A4A+38fG=85>Ve4<]HR=KCg[dU]be[>85Q1ZS41..aD1c&HU)B1X)/(CfbA=F(K
&\<W^A>3Me-6dP:CJ>_YOS6-?Peg)gbNEX3=:20eU8UCO;3\POF7B3PaT?AVPB\.
Q0H[4)]Q@J(?6E<^Yc&TUg=RG@&+Yb,DN.X:gO<)3_1.S5OaJKA]98aPZI#D+YM7
.X8]F6PJ#/PHYTZ6GJg6GL&0.,\.:8Q:P@TF_M,4A>7O#@IZUY,BJK3&6U/P_+AH
\:F,7PUZMRBgM0BR<9aRd-Q_Y#g#@Kg,R:V+9Fg3+]^T&F;NEWc]TO2[ca+EU@#3
8.UPQGbO9K;:a5[-,7JYP-gg&W_Q-PI75NB39U:4RX2P@M[cZa?\G<fRAZRgfMRc
#V<SbGU9DcZ[MP&Yb8e;&??D,Oa,:g2]R9#YR\aDCgKZW9QL-.0SA4.Y#KW7aA+&
:>Ib4]Uc#B^#73>CCe.S/C^DId0dJ<?Z[((P,<U@2L54=RZ92Z9JJ/::)E14ZD(9
IPUG5d234Kg+J8[Wa7<.(e0aL/D6J,?L\_ZSHJHK3cX4Z3?@-ec?LF41\;Q<&8TH
DbS)XTQTRa6N[]_L3FVO=1GLT.J&;),Wa?R_FHN=0:T[[/SX_-_M&C3?N12EQc2W
bf&&5JGM;N]C[DX:S;O^((gP7:;5QHa(1]R-)_-?OR=NB4=7KHNa\/J:&Sg(/5Sf
RR3<=,;QO>QEffCRG1E]/GU\gLYY8G:@1\3<&E,TP,FWPa8Q@YQJ8X8KO5(cAR43
#J8&6,2LdAdN;2UE6=94V^WP\]698^00_:0A)1VM/Z#N;_9+(3AcAJ5L7S0bJ8<A
UcIGd1911S2D0SBcJ2Z9]/GD5e:M6PD.\T5e\YP<8@/cP(X8b:aL\<2RaX3=60WS
GG5NU3BcXY?dAW:[cO9@)U)6f2/a#TXVg<?a,P_7:;\IM7_]^Df>c.OT)FJ>G06P
]&ED0[K)(gN<F\7Ie.34WM7+Q.YgLS&PKANWC)\g)(6W+d]NYK0I6TO#>,Ra9THg
1?44ZEcS>XT#]5WO4HZMR40KWT\a>6&96&0\YS38>4IQ-M,6T<(DbfD1&d8>D)_R
/>JIUE(W<;C3Q=e4aQ]TD&)R6UcVU(=2O?&KGVRa/G0[WEacQFTYH5c]Kg^29^HJ
M=[^),7;[+BFf&AO6b(E]WVL=.+F1ZCJY3SPY=FJ-6K:eW5+-2HHQTK0NfU2-Z<S
:1.E4@M5?YV@>U#5T/1?&]cR.Ua71W]_,H&9@>dA#JafQ=JW+#/-5L&,T09P)_1O
@Q=WTST-\E1dQ?NOF1BA,D_T4AP]b54_Ga@+NaGZB9J370H5E2\Ne6YR)+<TJCg5
?\INR.;,FNTSP^,<BDfY?R1#JPP,D7fD8Z#B#Y-;R><@GI9a9STg2GT<V7ZAHLDK
#A#f5SX&#fI=.Z9JMCQb(0]0VX;??LW6CO1c02N)^EGL]fE2E>H:1WA(REB=6D,9
K@0&JL<F=+PK14I9?eCRCD#dO71+N/ec,-+cK>,E4fdDXV]U\)A43&:>aS8##\N5
?G:c8X1L\:9f/#V2_<?/_RC+YL,FHIZ[cQf9GYBT)WMS<;@C[c5GS[TO^3;V<Z4V
V:@^#+:^Nd0H@9GO62XU#-g3]1ZN.HcZ,@]/W^_R>#=TC88AMN]Od0fWH]_P6L7@
bKB:5=BZcbCB,-^Y7M(3gHcJGU5Y>-;1e@<<J[FQ:T/6I#3JSPP-]YU6A^GfZ,cS
_9[6#@]g;Q[\L5,V6V1OLN4NR>9H&3fQS-e4@fQ>I/E<-]1;HL30FKVeN?>)^KSX
4>6S&VeO-:#D.>CEDYbe,3OACIEQN^Z6MMZHIRFHDX2\CTW@9;aHf#Adf<,b)f4g
dKVZe6d&69K\BIXBC.XP+N4K.Q:Ge7-bgPO:#FH0OQNZ2PAGQ7&F0VP,5LLF_YcX
J(P5.2_@CRMGP.=FB;38;c7>BHAQ;d\<.7#.D6f7&8MX[L@/g5W\a)Pb,\6f)K:J
\)(O?4ffD>4,^@W6&3e2a2[0(aQEaNV+U=DZ?R.ac5.f0-94?[HUfMQNP4FHL8KQ
Q]8M.c00ZQOgTKcYOE>QOK_d:(^)BVc3VZL30]XT#8;?V5/U-8fGW06Q50O)U=b.
Z(f-F3]?JMZUL>_A.2K^I,AE]8YHeeddLMGP#SYE+Uc(],F;X=6GS;N8E4;L>NC\
;CGbMD49c.#9_[:4<,(\W(>VO&;]M8UHB5(ePNY+?0[#N]Hg-X/9]?b8#;OcT)\#
+Z5.E\.KH1RYOU0(LJC&WSEFA;7FCQ4S?(#J0,+5aK6[O:N\Cc?0YD,=W2d:ED59
dU@K7WCS1AL<d>7<,4dV3-L(fNLD;)d#^(WMD)W9X=&QbI10@IZ3\ANKWG.g>bVW
KZ9..QXRDCHDgI:&2P-<:W;=eBN.[;/16N/-ZM&b(cJ6YE=.0&:/8GC=Jg@Z_@Fe
@/N4]eQ[V7>Hf&B0F),XU#KBg<2R6&?&]Q11.HBQV9,_1+9Q<0R4=6.C3J^D.gd#
K;PZ@J,9=4f#/a5CWTJT&F]IAC7d[KZRB#\K?M>8\)&=C,cGeT(ddL/Q>fD81-Od
&==A.Z2+SbXNaJ:Q+VgQ9V&[A8YG[ZP^^CG.c[[1V(P?QZVW4_8LUKH#QZ5)/RH>
dH=#9V\)]OC+<fK-8M:^Jb:&3YVYeNa&&eG/,KQULL#[Pd&^7f,-AP3BA]]@bHV>
8K?VCa\6&>[2[OW=3LH.e(W.[6QE8LT:;6/>ES2eEVCf]1>;ZNKE[Z3&?\GE9ZL)
M_>>,HCS94M4Z?NfJ6ZKDZL>XZA9fAGg5&Y2P:4bJ^NLT=C,/_W3^N3^ZBc]2da^
HMSVF;6^G]52gg?+6XISRc@.)eQDEg.V&.5(>_[][VTgX9GJS36:.,^N1&&#[_]?
R0^V>+\^+;EfW1XSAX#Uc7YBYZ,VSUH0GV&CGgOV,M<d<P8/RTD=<2W&DO4e0Ob6
U3:5b-/+DL3Y@TG?N&H+MX_ZQE4c<=.#<7/4?=F_fUT0C&Z19^+KYe4D9Y^&V/&Q
OgH8K#5P?7AU]2[>A8Bc(P+HCR[7HVE3eC2FX.01a@=U)@V3.3B]W2Q&54H]T=<d
7025QWbEII(C]1CLWES?bAO^Eg-b.X1X0J>HD\^OdXF0M57>^ZXB\:Hc#ZF^C?]V
GRPBO,UCYa20G)4Ye?HB&Tb=)Ua#3bLMg.^\W_;fW6;&a\I_gV16>[@N:VJV>#,.
.Y^S86B-.8]0E>H:BgAe(1GZGN7G0cRWM)b94XZE79X5ZU_C9cJ3/5YJ8]6;RdfN
MFdEe]FO[]=b,_494SBHH+bdHMf;]+6,/NCYV3_c>6_4AK8)dR]_9f:2?X;:/>8?
XSZA-LY@fW^DY.9&3EJY>Y:g__&;9:BEXg:M=(S=UN&bA#,;AYffG_U]M:8J7L0Z
e>S5K7#>[C<3CIKR4>a:T(NEb]60&E/,&R>U\0&dB:aWe+J(1,N>>Z<?C5U8KcdT
K3NBM^5Qg][?213H1S_gW6FSBX+D4?5;^&4BWSgXcDeb.KdSG)<M]8RNCM^UV,.d
0MX:(N=Q?4VXX)<;F7@C>0@fV-0NeQ:3^E,d7Y;Eaf7=\?3ZLH.[K=-G;6VG\>2G
<^Z?1.SD3=JIHULQ0b^>4O3dZ?^OQ7KO[7C-9ELG/>-?#3:C29g\+];2a2Eg.UHg
9XaN90d.3MNZG[N8S7&6Fb50MbQT7<#HS_ZTOD9\(>B2b.9C3.KK=TQ\=>H,P;H>
5Q)ZW=&HS98]CJTbPgQRe@,74?4)F.)U4bD#\02DCKQ=:a0]/]HW+O1?(A0f[DS1
FC9H13gBH205Y.:f\;;55W^)O3?Ed61c1XagMe+aLV=dQI,+^]P\@fZM#K-N9#WS
acLg_Pd;ZA]]];YSD0?V4->GJX/\d@(5XY)8Z.V_[)6I#G_.B.2[HISIGXA)(a:B
DCMFT7(ZA^A:0HT<.J+N.B+ZJZ@JO&XAbJ#K5),MNE@PQ/_)N])MLF:K0XD3@\Q+
QV[eMJ6S9O-;L]UHE&S;fW^HHYW8[cH=)TH[A]<cHP(O]-@&#d9<UPPJYD_CGS#R
/\N_805Ab;3=/,])28P(^<[GD</.O40[dgS]dgTeB7M[]3AdCg?55XO8+\+7@V@3
(XDL09P[CWI3TY@>NHT:P]A+W5B9=)?P)6-:BG;5g^Y:4[<4bD13;SH(E#&/e&P@
VAf/fO(E::?,HC^cf(gZWRZb#38=_DT>88Hc[eZ-8cEX,1P[XWROF4C2)=A)-3UT
5\YV:6IaMOdFU(#L+&XXC5DP(&D.FC)L7M^<([^7A+\GL&,\#[O>-^_I<L_)c:Q7
bI^RXJb8?B^.<]=J:.AJ/J,F)Y@IM-XNAX3L(ReQ?GWa)R;K4>8D_G&Z5[)AW5Zg
A_^KTbK5M/1J\3aHU3Yc4SC1:KaW(G6\\<S2feWJSPYg;HT[+gDZaMZ#^Bc>EG3I
U&R3aYX>X]CR[/#=)(g(ED^@c8g;aP<gKgg6TSGX2J&M\2(+bPWV&I8O1K:+Z2Mc
c=R&Z->[3g4>LF@)[c5\9299Db31MX?@_,_H&F_5?1I++TgbFE1149,T]E)<8&S@
BPF(R?1dB]\M(S+2c&R(K:=&I?5ZPLD8+c((b6E;KT]Dd.E_fNW+[I7)ZK6-c;Oa
5N_@?b^[ZTPL4\0-#Fe;#aM#&J;_4#_e&1g+7>,HHYOQJb0,@,G^R[GQ5#b6096(
Cc@G-#OOeK6KR[.FI(.;\8_JB]0^?PIYe?#HJ[PC[<C>M3TA&;:BG;RfQP(dOgBF
b[\BLESNKR;ANYYa8R.2QKTf,2++.gAI;S_A7eH(6CK^G6K?;\-WLE?871RB-4-P
GcPVUK9J)S)+-DX4C>.R7SHOW&0=X>AI\[0G6&TLCeU:,;HRe6JfRYJ_<Bb3O&OL
FSZ[./S(P@a2U^SUV<<A36fB\WaNH8E+\A5.67P[B#XOU+e\>a2#(Z(eROE<]HX<
XV[;](^@Bf_<b;\C\OB^5HX@;HZ3QAFV#03KU:70\OE0+.O9\98D\KBP(?S/=T3_
4;W\<<gBIE#KCN#NGI,]bVG9B3/6G_eXAL#0_DUZ0\-,X=Q&8VX\H<eS?T)P(MA=
Q[G=Qa>(XZG+db/D\L&_KVeX<,78WWC6[-0IO->9<:MFQa7.c0Hag9K=aPAEcF4X
OR4DP_eS6K;/+QXP2)853N:<g1Q\Z>\79@S9<^Z24BJb@V^f+<#IT9(&R)L(O6/@
/-4^J9X387F(E;Mc9aR;PRc37_SEI_#A;]PB/>).#1F?Xf6VK@#YP^d1#YP?c,45
eGe[&(8I1FJQY)FJS1MbTX++UEIG]IHX5?E:-?]53YX^2\VMDFLS>&_.Y@.)Z6/W
(D0&MJ-#WZ8Z[MOWX;K.N#XI/SF9C(7KEA<N9T&7g;4[OGQI2H8^bf@/R0[=@^ZZ
2Z#bDOE8S;D6@NRMXUdb9FB6P0^J&.Q+Z(0+<@Z)T(8\fKT^=E()b(GH#=9fUR1X
b_WP1T@cAYf\-=_@8LP)JcIgLba=A-=T80,GYMBW@ALGE5HNIO?<EDfDK#H\KI=>
c@0,5DM@DD42L\.JSd+_V-;c.J5^Xg>-5#:)#XJOCL#]AVZ3NHIN/AS1dTOPPd<;
J[D)Q1ZJR2,:&3f+eW:A;ER>f1_K42=2^NDcXd(\C:g=b0@2Y84Ga6KQ>SRX6^T4
).Ie,8c^FbXG6>RA[>3>F5P0W.cI\GgOb5ZQT<9/&+IK]-^?Z>NO0/F)XQgcf2(R
@eJc>?Xd=#,cX@RO(dKS:LF#fOUT^5Lfe8@@bQMDd2aVCMKGVUI(L<\9Q\dX?:-Z
IU;/AdQg)YB7a,E@OL9P3T.eVK1L@Yac9ISY27PM[2T@\.+^)=?:5C6(1e6=8W,G
UMff:Q=C(aKWTY)a6Tg7Fg3c]K-3;V^0Vg]Gf4,T_+M+B_[[?[&c?P?=)^RH:YN(
9C5S/S@VcO=&6TT25d=[BE;GQH@-C,X2NOI4,Z9C09<7>/(8:LZ,-_,1a(]^F)AL
OI_b9+O(2&[D0JbI7f,I&-O[g@WUXLJ_;FBLGBDe;>MB.4/]_geW+Ve-K^WRZN1,
?1.6dN[.>WU)HM@a8VPGcBX]QO^T/B+/B3VD&6f^dJ<>K7VVfJH):#5A?W97+/ML
)6U6=0fH5J=,5LHU[SE07.X3W;VMAd#8C#C(B<B+#M32Q13.EC8[1Y2]?VW08bVE
HC<1/OW;J^MD5\e08/:^?5:=GKLK#EfE<QV</<#61Hf(UgNKLR0-D#KFG@M_GPLZ
bM/3>GfA(6C+QYJ.5c@DQ.E,f)K_ccN)gZO.OX-[>GNB#0UT/cS/H;9gH]UT3I)3
SDBI7-03Zc_gAMUD.f;a\a>3ZU4S>[)N_V,&>CFe?F6LXY0-(MU<_FWR43B\\]D:
g^XVG_^?1=@@32BPVMXH+.(Z3dM;H,eY,,80@+J:G\9\X6V<75R[:.H(9447S9[[
fU9[AE1W<_BK6]2Lc#G,_L2ggR5#3U^)Q.LKWOC\eQ6cQG0CXdMK-55RW_?>bK&(
3,TFOL\PgB2C5O0=-S97)XN6QK4b.Y\AfQK^05eRZ=a6C<G/S0JS</:)>WVdJXXd
_,:O7X&T:;H9HCgWZ(>(H#LHD0Ab+<RGX9+\B8_dWUZ.7OA7fN\DXYZOFH0R?>T,
EL73B<U@61#5)+>T^YS5++VSeNGa?/:L.3B:@;>1OXR5c:LXf+X4bY;&(?AQ>>(#
&,[,JQaO9ES6Q6Q5L+[S6]+VZ7PPC/1f[Ug@Hf4d8T9I8@ZP2d[3d1BF3_c.:/[G
e@G+)08D;d[IUY4WfT^<?9bV+I9_Q]\0_bDNFFE4b(F575HeMQ4SI=\6K6)C_4:=
3d<.4#MY\M>(VHLD0<EZbaSFO8Ve;_]E?)Ve6TDR)_/C]T17caAg72SV@?(fM],3
C?USW/H1+>X2I#,EA6QTc#(W)O&Ec.a6bK3\-P_?W77[;MH@C)A[7BFB(.\08)[\
WZ_L5)1YB>H>bSFad/-R+:Z3e1AZ<OM74,5IdA?TEKNcIf]B0?=A&8UGF2bZcGZV
\+2dUR+KQE\W;M</IfM:.4//:5K<])K4<][Jbf-GPKB?f@RU;N7GSA0NA.O74F8W
CZe5BaSg,3:4fJ4&#CD-PQRa@SdZOY&OFb::eY?@VSCQ)M[R8FQ95W=NC;8-(I4/
U5L78D1I2fac:5&7@O9@Oa8.<5Ze>Y]I=[Oe?RTT6>-37VE,\1+BR,&)TKYOP(H8
WQO[NcJNN(dbC9M8;QJ&eNW;B\D_=UbYBUcUE1#&#._6>.K+BGJYaYWEHK;:-BVH
XR638D;eC4MG9]@RMEcPHD[3@E3TWU:T3L<;ZeMODf@(HcXH7geT(7\VCI:bOJ45
GXTba5-SI[5;LGXO-d,=RC^abOb=9<Q_D7UeA6,W4a-+bdI.bR<U>L<eRW/HQ.Pc
gCANLC\.95O>Xg[71b8H_6ZGaC(3MKKF61e_[A]A-[VE_,N9,\J<KJ]0N<\a.3([
7S4735dW13OJDI+7Id^S@b9SX]JaOIV0D:W-)_3;-T@RI+^8O?RdOd78=E/K:e8@
;9?C?#XCZIO@U/OB=K&7aXVd;J6fZB;a:8WHLCU=?fIe,2&PdCSfPX6I^SO_?&6A
86WIRUA)MF))2H.K>HO8Y>bAG88R\U-P=:1A;AAgR<Q>=N3.)(77YP.CI]7L]/ZR
KXed=fb\d1+#/C.1#.#dRO^c9aPQ-VF<#KBc4YdgWD=FMB+G5O>H/JW7DHd987L9
]PJbf)1P3]QYW?30I8KQFa<I]YXE_9.Y3^f9XGIc0D^P6d9-##MOG0RVH2Q+>U4a
DZ10+P]_P+1;a(g?-\B63+SYc8eYDcH:+MN[5/1,aeaD=RR+6NI2A7(JaS(77875
KAf;de0XFCE?^f^_-8/Z]#;R0[;J-&>(_QA0d/G=1If7HEGAa:CKdV=@FafGMB5B
bRgWd<5_;?S9a>>EN9E\<UZADUJd&FOAD(L==CK[P7DRK<4;/aSD@UAJ@6H]J0J=
KS^A.(UVN=8C=ZW/Pc=Z5^SM^I(FMJ79cIPH6>Sd-]S[C#ZPS\N[ef)(S>P(S=T5
H6gK?:M;U42-UaF=+W+T)37MH55\L.1ZTUdM:c>/:R(CS,CXLM7)#D.gW)Q>8X[@
db5B(4XNH&H:/7K[UW8AfeAOg[(S=S4[+XQ#RUD,QVFT@:Y1Q/d#PeY/B4C8-=[]
a-K\<(/<\WN(ac:8-B5b5#@=WH9BJ0f=L#H0Lb-:7a,cK31+LQ4\<9RF+FLW;]B4
Q#ZYT5?dafRK4[+PDeG1e/aOQeCN=93Hb7b)I,RNO^>^A3cIMXY\8ZM-NPV7^NZE
V&c/a.\=_Cd](0MXf;XF/OMc>2;b295ObW,46dBg-3G;XDRCW,L6[:X84\\8:6d2
Mf_-4>V<I<Z(<)SB?GZK>B:^E/G5S8\Qf@Icf-HC0V<MSTB+K&4L9)C>O<:19TIc
BI@=F7N;L+EZb)70>a1M9J)FRK)2^g4C1\WYg;gZZ1W5JN;eIN9O?gJY=VeWY@@<
d&C7Oa;P^KPbKdN8gZY5^4fEZKV./AWI=AbU;VRe>,#.5L=MB)<S5X.cga;>2I]Z
:744I2>5Gg[2.beTgeeDd:)a4S)gde)=SAU0;^[GYLYP#G<NS,-_g+^X&Q(f&WCb
8AY0e.VEFd#T3(7:/(GSF\a=MI@=O6T[e)R(ZNL5<&S(HeV]ARX-c?@.;<+B)NTD
Y\C3Z0<a3G.#[LgA^gH^:>EXS2<7)]^VEV^U:f:+W))9<;-2HgB;7&]OXU0YK8NT
gJ94dF=Gf-ZHKJ<>>FFVN,IRJ[/(bdg.;_H:SaW/>1CMLHfWE_agX3<F\WVJCfGe
9^Y>Ua;8QMG7O>cd>E8PW@IP[=+SZQ=-Ee8_<e&D+?IEH\0E-\91SVBa#-74[K<d
d]]P^ef?FVS540N=/-:5E&BWeg_H#g_WL7aE&=fG\7.5;[E)DV;;@C]:VIfP)&2g
]T9ZCIC]>b0EPbE,K1&..@#SE4aE3K0-VNZ^+<72edO&^^#\M)&@U/\[P:ALI^LA
CcQF>9,M]2b)]P7@,2Z1NdKBR?I0Nb.N^KH:42PH54(]5+EL[B7L82gaZP//AU/?
_;J=8JaOd/EOCPMNC15_-:7/T5:NK&a?P>YS-IK,VJA&Kb6LdM(@@cYg>/T7O^IQ
+9=UA==X5cN7X),;.SMa7<UN:9K7W0SBXQMaW#++S^\\R_E01]/UcD158dE.3MU]
E+W0]9NRW2UT2YaEUcX\&d1AW-cMEP<<JV\;00@PG?PN&?_]1>g/>^\JWS&J&QO_
US@L1cRV9S1R<d&2Q>;,HYLM^La[AWS,7/I;Y?e1f^+>K3e=Z&<Y&T43UMR.GD;9
?gF]BNJg4.DBf4M_PM2SZ\:cMA][cUIATY5ZO-KV-SM^I-Q2g1<f/8BYSd@L4V1P
P+G6O0Sd+caaSd2=0A/@D4Hc38d1:(YRT8EG]30##e^2<NR3=N3@e#cI3aaZS@]Y
__A&#4P?/8^=V:HaZ#>F19@cN3RQ86QE^<8CT,D5a#FQ/@J:[_^TA^CU<c[OB[F<
/.VP@UXF2BRMC@0dIVe^6(:3f4Df)]c>.)DG<=3\Gd/F#dW@+g&;4ZRLPAP-K=KQ
\;;Z?APgG=/I6D;RQ5f[D.R.Y9.[>HMUeJ)3.HB9Kb-a1Z.L7#W6<.C7QCOTSO^9
)_UR;F7VZN345WT&/&#Q50b4ZcJa2J,IK4KfIOHIM)Dc4H#9NRACG6;ZCWe=Cd4]
cV]VC[YITG/-RM6@(F1^GR8>F^ZGWE-]-/\X3Q=P.aQD=fA=0gHD?AF;OA\B/Od3
R/9g,O@FU]3>.ND&M7MRT2Q@OSU0VcZ1,YKO;+_=W,a_0K\-3]@g::J7E#GI^&)g
7.XJJXQDA>)Q:;714ZbdP1-=/<XM>@R5NA4H.cc_W/<3VT=A(:5BY(269FRdG;NF
S?B[E.aLLS_=a)@/YLE:8=KaYC44d-&NOFDUZ/X[S,:fgR^80ZbFfeWI1P@:[BZK
ZW^DZW.:425W2\BFOO?,J7V2e&Id8_T#Y8&P(:aNW@aE:ad5PSQV1\FQ4?LD<<@@
c=<Ud\3\dA[G<g7N3#:RZ60OMWG#C_<JgW5K=d];@d<1&#?:Z^4e39<L#XeDdTN]
7MBgCX<f@-8=5&1+@PML\FE2?#8SKPeM9;;8.L.,bW?T(.<X7JIY7G:Mc;/B/CW[
DGT#)-UU?f^QYebdKZ,2M)1:aO-3XACMg:N+0KL>C^+E[9I?<H)X]Ga[X0JfFAga
80d9+F]Yf18P[UV\&VP+OP23(3E,8)0?W2>Q_>5fLQ/V/XAJD/VJ0NL&37@.T<+&
42?Ee]>OB2BG>0FP_)IX+,\QEcZd@ZR2c3R^V(SIef[?P=GQH50H\^6V2.L+XNE=
Y)RO75ffC.]N,dML<F>TR:b(#C::^3JB9Jb0\H/aG9\g,_^(5RNfga3YZ7CBEH,Q
>,)XI?]f#SNYSH@@W>@SEZeT--Ze@WBC8.+d9EEeFT0\@B=#<1?9JT8AZM>S1M4[
5OZ_W4B+7a:Z)HcDIO03XJ)U#?DHOY1H+2<9,=F/?_6D,ZCLaHRODUWF6c&07)H+
7e0<RNZX@0H<U&/4.IdRW10K/;K(KK_DVf(-8,BOQV:P7,R_9=:6fE43.M_E[X[C
(1[4&DZ-ef;DN2,.2CN1@E/c_2<Bb=-Pd?2)6Ma(B.CQZCdE-]Ve6\3cK?#/S.S)
3gQ)J?8a1:3d>6-9P\HFb.(5T0\M6]HV)Z@bJE[e.GH1U3d3bdP821O^O4LN0T[A
9D\5S7^C?b_L/OC=K&KZ9JB-4&g0UW5<gS?1F;EY1&:bUd;;2JD_5aT[S</N9.T;
W])G79bY]Hg0IGS-Af/fV5@NGK+=AE/=Q0Hc(>8b[?4UU5AOKD3H.TOIdDg(X3:J
b[^OdY:B2P1,=cYYbLPCEEP=G.W,@W1)P:])(1HC=TAgKXCSgYRLEIFcX+.]Lb][
HgG_U1(2.ZbW0OWT7AR>UWG,=WQ>e1#bIQeB@0U[J@\GYVN8PO+30>G#e#WO2XJ.
\ECHT&[SaOIL/TdM?Z6NBWDZD2SOb^CC^HC]&JF=P]#]_Feb+Z<1Z+1()^UZ5#W\
.d:UW5.S^)dAD@b9Y\DKb93O#;:KROTL68d_?7)_S=)S(Db>Jf<PL^OX]&>IVb-a
O2L1Y?ITVVe,7g=H3.WCXZ\D@T>)P/UF=C:]]/OX0g/#,d])ad61c(_UJY+ENeO9
Q,?45]RR1R#5]X]?XK]GEPE+(^><W2abYUJD&9c^BUM6\d8(@QVf3->8Oa=^S/\#
;;T9RCPeXbMHbZX59#e4EYDa@>?2>@(O+;G>-C7VW8ONg>JQFHEdY?MPK_91f3=9
@^O_f:U5TKNSZ5B-b([bE+>Tce.Ma[^FNgdYFE[L6@\.VOC7^P0LPBM6dZcU(?;9
G1B16E0P/Y^d^E1_V)]c59;OLJZU9eBdNRF3Z;].?BXfHVKFX^,#JP9ePIDITYaK
T70fWHDW>-@GQNfIKT#8^N?/AO(T0)JF5)3Zac+YDWZOGSV4PWU\:ORFR-^2^0O7
9GJ@NLQ3=WKHXg\L3XBAW74)5&F]#3^S#ARea;\_50Z;E,(+8>Q-&>9C8=8^DDP]
.a02N0f6Edgb+K:9(3b>DAQ:/50I<B_\XWcb74>g&EC(8+NgXSG:BDLHI[U98)2O
NG<3-CbJ=@IUNd)IFg_JN,5.Ua5K]T:88ZAC05@eBcdQRNTeM/9LU-:bJIPBS+MW
ZS]K:8N-YN8]_J&cV]-56--]&a0X_W?]B77XdHS#9@#).f1?I.TRW38\9;AZX0^D
O7BbR815KY&T)TV,;8MSYbFQRL<F95gO#:8YK?_DJ.B+8]Q/C8fYb1QC^Pa];AH<
X1c6.PU#WZaEC4bBR?U^B#[ADb^S2A7A;K7O]0V-7a5)EZX:P0ZG9,@/O:?EcH1D
[HEa+/(@59>W6BTRCKHOV2\+TdORR\=^Of4UbW_O(b2b:K.aA0#c^P7U1U;dQ\=9
7]_A;RfU6>R1@:0-dN?/Q4F>0-VMKeCeZC<JKI04#\JZ)Q1dgQU#aZZZZ]]P2bB>
cT6bJ]0).Uc_]fgbU.e?#Y);DUGG.8<LdeD>3>#^f<g3S[W5#A=Q8PV1K-]ePQTB
:e#58cY6AFO_^Y4J.O0d/1H\fMF3P<a#Uf&?T(H@b.[J^0(BEKg<<fGAgZ@A39dM
C5U4)e6SYIgF>7G&XBaLCf_/>?29Ib#L30GfL6L(?S\SAV<\90G7Yg8A_?4AFRdD
DGWceQb5T)<CdS@fI:\[ADH)HNQ<^@F-gE64Sg,J?^S0U[P&H(&gB>HA])AH+AZZ
K?.QZ3[[,PcN;-X;P;8GbDRJ..M1-C95I=?K_#I;4C-;I^YCN8:0/_:>W]H.V0W2
b=.LGURX#d/03E+PGL9bMM;AT-fHCb#f?.40K76NE+^#0,XU)gd@fX-JFWG^g1&^
9b03e#F^+g[+7QW@9^_,S.1gc>AEB5g_;/5cG6PEONV07@;A2.9A@#=JLO#<L8=/
=I9f+#AfKJc#6L)47-IE+bT\f[(b&OD0]M/e71D)EePENBa@7R1#A,:YEF<0ZL+:
3=Y)@W2gO,ID9=G7)R&\+YCeM_[_BWN?gJ384N@YVY&I#cFYQL(2a7B5fQ6ObAI_
FRO&?JQV66TeTbgGZ?5&g5HX;Q(FJVLY6<07NB@^X_3QGA609T96Y90Y5)VG\MSa
PRI,0./LPTOOCYVG@,FGC-@UJZB-]dZ\(_\;(H^9;INB7U8d\R?.1ZE.D9/F<a08
3Da],@A8@2I3^]5L;8.)[#6E@JIY/S/#8^XW>MR;UXBK#-(O3(+4W?]B?_+A1bLC
S3,Y<#fFdK<A<&-L@&#cfXaJYC)4,GVDR0QUQg5SJ:129fW(T5=(eHeZIA0B+a.?
\Q=W3(^5U;BCZb@[@Fee=@_8d6^^^c=EH@JV)A0)@QC[fdB70/a/B2ASN)>1D[B7
IAL<b^L_4?HWKQY>+3=eA95EaW;b,_<DFGDNI(V,_1@YaG0fG=+0<E)5>A+P/(@1
1-21Z;2@^TD?Kf_@V)\9Lf>OCUMUTaB+J(.N2fgc.SBdc_>635MD@(D]N^=,>d4,
TYFX7^#B20?/S<;\\5_RdTRM1TSfe+<gO.(/-H(UF.R4DNV-=Sf--.5#T>.(M<Q7
N.\&cAY(T-7e8_?:D_,LLLVEe=dX#\8PH-0<gT;UBVQa\.NOOcWRPS20=,N;LTQW
O7E)d569M_D\g06FLe9aR1SW8V?IQL-SVH8E75/=MC(9XRRP7^.9R+I4f^UR9#2R
)Y^+/E&^,[P4Ac?M6>Y(]A>E61[<9>/_:ER[UX)IT)O8.5L0EK(FRg/2&FfdZOU\
^PcPR=;\#^bYbMZ<c0+:GEd63Q]Y>>]fd8Q+_;H62901E(d_T-+EJ)+?[D7+I@0[
L;;BD:U&9_A^C=Bg9f7-<S0dZ,(5R0g]\?ISCYXEJdG4,46-VW9O6PH@[PS3B<?4
30I3SA2MA+\)Bb=db]/QO@H7>P;),#_M(&05KQWFJC:>c;<d7TCCP8X<,V#6JPe7
98aSN;DZ#XGE3(H)7>&1\VXM\Nc4g[3I[P\VXfc1#XdK9CRb1@-aQBI9Y^BJg16:
F7W;VTf8Zg;_[CH6Q[U(,BgV??17@aaL9W/)4NQKWb0dFSeKB:fYHE2YY&EJ_c=B
Yf:]7.624DY?9,T=)6_IV,b?:MU]1N3[-L9aeR^.10.9=8N.>^7;)DYL1OeefY4N
-WSJ<G^.O48:e+<aLP=)Z:@g(]QPE6aa9UZU2>BWDO&?B:)VbV7HU>8[\\6-M)^<
_C>H>#5C;8S1.M<YR3\QVH7-&25_.-:SFF_9\.P3a4_@90b2fV2QgE/1=HHaQ^ZZ
fOG5e[QJA+HVEbeg:YX(.,Jg>KYHREcaK8F(B)UF>7NB-WS\9Q5SdUX<fRZ57Z#Q
BJHFTPUeAFV7._MTGgL#84P:=4FRd/47B&F00L]6Zb.I0:LX;6.bd]82)gM85D#F
/P;,<W5W&<YJ057PXG^P@eJ.cf:&XV)]&<\FPbH?d=Cb]4?VP)H(;4>975N]=HA3
Q2:B6:5Y[-A4HLTPUHdK\NVP@.#:cfgEBCT@:/dH9:W;DM^7\4C65;.SCVDZ.\@S
RF5/-H#YRHRd__GB24YUcZd-CMbcafW3V@1-D^I_0(JGa-GUT]dQAfbL+Z5,Ac/W
O@>cXd#Ue1SF(3Z-Q3ECFYU9VE0Z\.XfV8.E[,5Q8eCV7\>eWD:@NH[FOUN:Z29_
2[Z,e0K8XDc=CgU<1]22NI295H6dPQaK>]^LWc(AbTN#FeX9_//5L_gJ32gMIbS)
+M>/>Z2/EE9KK.7K3K>YW&+.^f8N5,b(9eK>MAB;5\T8Ab8D,]f:8&\_J?R^YEDH
2V28Cf33V:Y./E-Z<aNG8;J99#acDCB^5G4d<,Z^\@=/@gfLgM^3?-#R;,C=\Ge1
#aF6^(gH))[Zf^DIbJV,E?7(RSRPVUe)a09K]aG#_&Ye1d)]Y>B2bETIA?+;>@=4
a]Jee,OcWfS\#8S;F2[9@:^g&0@>P@0=@@YGbJ5]@NXW<5UVNR=D@Wf.>@F1gONC
/_2_3>1E?WGG<TEWb?3F;Q>E#Mc@+&ULfJHS7e):1PHD\]]J6\?U+U<[=ITPUL[J
)F\;8VOT[C2gYJa3?N-a&d8^S8^C7IDfE.d1Ngb#M^(47@R9I(,U/#Y12D\(Q&]>
RP<L5.Y36B]6W8<WCWL(E.K.V;6OH0L>RD6.&.CR(YC/Q@HDJN5b2D1-9]PWI7gC
>(:IgGB3PK9;Pa-BTdM_/)ZF]+;W\@1&3gU)/]A]FCR[,A6V4J:=27+I_8:2SG.G
D]?LSEU@D^,9X^(_T=MPQO49N>6KPQ<M^Y?CaQ;<M=M_U&3Y6=K&e1/@&;=L\A2K
0cMD#)BLR>LS0d\O:R1L=QRd3Nf52OQ>#,ZEEX:J3ZQY(D<5LS5KS771^N24KY\&
S(8JcbJg2?T#Y_AE_(GZ=-S/+0:+Q74STO7_^<YT31e<4Y&\La]L@<#^:V/,YO3+
PR#))C-M2N.8T3)2U@CDO3AQe#[_/OF+W/6N#^<^b3Y.TQBaF<XC#0@0g>e=9SK(
(DeUHf-aD:.RLE5\^5KUH:;UMU0V78O+R]dJN[3Q\)LFD10.WE_8-\\a#[e)CAFI
V2]/2:9CE/>G_W)U&M(M:=?>?-D54,PNISAL\VM,[#K-MCMSH1b=gV]g6:WdJA3M
6+EW:6@3]:.a28d7@E1>.L^RaN&cW5=TJ?#6TR-S#[NGe<?1e/b5-LZBJ+;/<&L<
,4ea?Qb[9_1-3K7c7M1,SJGc[?VBDHG3.G;NG-S[J2cM6>^9[]Z5f,)0M#AC.LK6
CbQ.TW[.P&/?gG#N8G^9fE\);94_;)V/<W^.NK,R1>JE0VDY:cG]e_8D?5XA3F#2
(W.d,0N66K7PaH-D1[.KQN=KM2=X^,,\+4&b>;^[ZP)KAQ-DLG\VACOeGc0WTA_#
bY0M[BC51>XW@)&1F0VX&68agMA>AIYU_@U@J-._]#V=,<Y5PIEe\Z)N8D(\OC\N
-4T(UX&K]>.M(FLVYX9\A@I+IOHaH-3/(C8\b^8._A4RK_@La)Kc?@73_1>Pa<E5
H,A5Y]PAKJM5ZY7HJ;DXA^<1M4J=:7XA7DD)SUJ?;T,-D+RNP77ZFNX9Tg,>/d7@
RY,<9PT)^cV@M1B709S\JE#RedFGO_@K)OM\<gc\4T?@g:f=-79OHRS)I\JG#7<;
SS-3V+N8\@#E7gZOHO4HB[d>V_877GQXEGaQJX&e<1-fOdI1CMB3U;EX[SL=,QM#
I44IM0Z)0eXC&YM;D5RU@6VK4gCHO.WA.C\)+??XI<;b(3=(S3/K8f,>0SECOgd+
V,DR_:(XTW2A0Tf_&\FgZb.UP>gcQD<L.1;A^+@AIK.A-9F4D/N&7Kd.g;=eARX)
YJIgVXMYM,Ye,c]gAYATT+2G@4V?5=J#,/&+M;<+REfL(-MPU01EMF1AS<NC\ebC
(]UG46Z<bU_WKV(J1IJ-Y00e4PU(?LEEVId7<KP@;b0UO6KW?f:]XXFd4.Cf]AcX
-._MaOFRa8dDLN9,2B0gg2[NR)2RBE6,5Qb7eIK7LYJ?Y.PFc+OIFU,0)(X.bTOH
[_.QXM49f>d6>^-#>Y=#&6#^Y-@&_cW-c=J4Xb1<[U^7DM&FJ-+;c??G,1EN7_Z,
W,(11=a0@R.<]UTX+AFF;#/AZT)fE/)UG3Y2V\I@9[BH=;UI20CY7;@]ZM/8&VX8
I/;&:C&H+CG-5>LGeN;4N/[-:KL?1A@5a3QPX>]DT(RHIALEC[C.d-e<P0O9I,DC
4P&f4HA#W[;DP<beI[&dX<;,RLV1/\b3>&57X9b:ML&VWO([+>51YQ=\<)4.ILGQ
@[-SOC]MPW_e:[.])bGI2H<gcXD(Zg59W?NYU\2RHZe/dMKV>I_aZJWPJZZ:UWLV
cb7V9/-.0OBId.(b871GZRG49ba]9YLa/Z41?R8V&3MW?CbPKOI2O<)W;Ie4@98-
EW-@PAgR7<b:3@6X./+d]VP5Ac8eSM+eV>+a,9SPA]:VVQgQM)B_1F-K\<fT[4XN
IJM0U4=E&@NB[[,ORaLHK79;1R7UbCdCUg[LE)?-LNXD7P#M?SIWSO]EK#dS#75#
LXKPK(eU?O3.WI0J7Rc5BP-^4Q0</L^[ULCKIYeQ;/NI]I&?+gY4.P?gI=^NZL\T
=Z@(V86eBK&PA7K)cJ\=M>2Ka17+M.V4@RLE;37JAL.3C7MJa1aUV8bc?B6V.#?X
>YH5-6_N<VJ\=U[LcXb]NSG;N0bc7;4G_cWLaL4)-V0g_.2c/SPX\EU:5#8CBP>4
36,?B\c+4JXe#]##WM]dH-8(HPURdbd957=V^K_4B=R2/]JNIa,JRGfY-8e\5\E6
^d<&[/HW\b9W&R(I^&@_HNM/Qb<P<PH1Q->&J(CC0NfB4.37D]_RA67I@I=U=4ZZ
(15\&g8N&R<1L_O[c-;/YcCDU@7#XE[;PEZO9Xc-AO>?:ZO\L3VIS0.\3CH5RVS]
T6TFT::0,E8_\0+e/_O3UY[be--I62AG/J=aUR:RcFU[2)&F1:f;eC[aUd;6.MLJ
UP2W_F6=8IWRZ7;XW]S1[N8>5Q&80=V_gG@FX++@;(PQTePK37@@UUL;OTSF1Pd0
]3JWJ#;(:>QDJ1YLO[PeI44-C81\:Jgb:(RE#aY_[),e=a]B6HL6F78&Z\<5J8Q1
Rf-)GSSEB6+#8+:2+TWf<XWL/(PQ(c+[SF>e4?05WKX_>VJ_O-/O>Ga0Y.D)#;Ag
6667=Z[Bd?50@H6I1:EPW4Cd_\BKC42JK9=Q.3cO3=7aAUbc^H1cOAe-BC<ae]]0
Q1-@S)L#/PVA6;MMRbI_7=/7^90CADe6N0QF,g05WBeLg]E=/Y@AWK+P]#RN9?_W
P9AD^MF2]M7Y.KD#.bQeK4&4I=4?L98^1NadJ(O-V^Sc^dWU9&\IHc=adZTEAI9R
\HC&9(Z/Ead09Eg963[F<c)R]>01QU.a7A<.+;WO\Og2Q_A_Z03;,&J^EK0fcCf)
3<^.f2e8(+VVO;I9b3KKSZ/9[;bb8a+UM>Y?&Jcc,-_ZEYPON0fNT:9bU/L^_ZH6
R/g[3Yd@N.6.M\?7_,<CGKR-JV.b/b?S5Oa@>D)dFJFNV)dCV7)UNeHIMS0C<a7A
ZPbAA417d1D+K34C+O0W.\5FY-dY9?2:FE_UJcfY?g<PY&Zd81XF_OZVIJ25=@P4
7PD#_A/]5IcM\,L<[T]PMZ6e^#9_8+X8^Z;bH,3/ZJ0?Q;FT.-LA=_OSB^DdU6V>
F+3e-Lg7=VNZV5b+088@B^0E9b:&PL[]T8e.?e[/Jg#,WJR7D_\eF)K4N+/[Og(8
+UYJ&;N.R(0.0ZDR\C)<KD,&63FY+-Q3\b?3P),X/;I>E?ff<AJ<OZ12ZbdKB+81
Je+@Ie^&IIFY(4DB[VFA+DRZ8DR,S=@b\8I2Y[ZB>#<S._N.\?)HY:C8KVUE4)1C
&>ODb0P7?+IKEDZ]^[20]G(geB2dM3=A]HfW-12V&3&CV_LLbdP13U2;<HS&dN5=
+:RB3;X,9>gEFQVd+V0HAQC[-U315J.cE8.;cVALII&=K6BQ\IL\WD(U4,IP6VeT
ZO]gQYZ3KPSEXgUPP/OcWF=gD#]8b2/bWe3X(_YP2&-::##9^Y6Acab[J\FS4EOc
25<SY[_5+@4Y#;_]TBaWQ4N:+KV96>#X=6J>BJ>cD#+#:KJfa765@<D)?25E5\YZ
3QEY52==:5c&3F&J-LK8YIU/[3(SZ<468\#,,1F\,ICc]0Zf/gH7]-AM5RNQYD>N
&fVaN/(3\9>+PS3GT>I6@E71(TQ]55_SUaK0O;I;Q3-b[DNN=@HLUe@=FM./R8^^
W-V.&5-#1G?8F.N6H,Nf5aZ+H>:);Y]eBfa@Ca;CC(g6D\A&((FOS?<(K4WH9-Z,
Q0g#+gI);J=>3]C=(QHdXc5Ta5Ub]aU3=6=@9?92>4daL9&=XY\U;EO_d,-X&Rd_
(\9+=5@VGS^dgU+UCWR[T4P_SP,W40D8e6U/dOQa-PbMQaWDU>(c6fMR+^7G76DW
fYH4H&V^F&8g3F6,M.3O5O2AL7>M#X#E1,R>UJ^K#\AKG>KU<L6<KO]ZUc@@P]gW
&-dHE7Mf9AKZB(+d;f;-6OScNCK:64VXK>gYBa3P/)8b^JXKP_H9@U&_OA6-G>3[
:b?Gd-.B_:UL<-@Z+T#HMb2aGI-#0N5R6/Le7Z?EUTB<P?NPE]X,ebQNb-d&Qc@6
A03Q;?CV]W_b&DMI:J3B@/[/:_V/52bVU_]:;Af<7@b>R&T[L_H-(faV#Y::DAB4
g2-&TdWTLedLI0+GU3R>gAeW,LRAI-f;7d]FJQdFgK>T]6Ue6L8.Q..+4WgRH9-/
@JC^\OO4?7[0QbP_S7V)aDcgGUEfdT0bBH1ER<gA-Td8<5#ICT3UI_V>N(5\?WH+
T:QD((7N.-C8)Y1=KD.;>+^D,=#4Cgd4W1ZV)AR58b6+:e:gAWdgQ3.22.OJCcC<
I+S9F-9GEN:BAfLKfN2LQJ#>>.aQPMSd^=>3Y0,Wc_]JKXNbA>ceVA?]F9YBHf(M
.bK,\L8FQ^L)5H-VJ97\/-d-_K-(GYC+L??+^R;D(@9Y3]4a4Y])I(RD[X+)aN.V
,O@ZXH]VLW4GEJIU_\\@Zb2(3LUD6D@RZ.(0+?9<IYE-^B?EQPD1Oc=]X#HYMX:3
(_1eb[,9O4EO][HC-2GFLJVNUGf)SN;2+#_GZ4@MDf;1FNcTJ#YP)8>Ve.E,YVSY
gLgV?6/dIZfWa[NEZ1b4)(#cFP^SGY#MDe(BWgPPPff^2?7TTSLTS=c+9(AY;,f[
#I4fbY^CbGEF.WICZJ=(+PC_[YMLde-;LZc5R4g7@U<,c_=I?_a^Q:@BEK08>a)P
e;DY[SY;#e;N364D,e5&)QSgfURWLU]LH^^M-(C6Of<I./9V;XKS;9:J:DXUJ.^g
:Q2FI5fRPc(UE[#SHA][WHZ@#g0FG\QF(^F4Of#aN+1V__=JBdd>QbD5<dP:U]VR
ccQ>Y>T33A\CX^aVJ&C+SMEF]I=/7&RZ)4NSTJ699e98cMA>/B2?P@N_0J,L\HQU
.A0U&H4O<YT[b7)X8]0B;:QGa\e6WXaK[B76gOLG2b2-KaEc;=(7BNe\f87J;X,B
8AE#NEaYXH4)L;F[]NQSTGNLN[Y6ag<+c:)<@HLbWJPTc@TE:EP/4TOH+U]KX#ZX
[55RfD[+2Y=Z5X35^9F1d>4L&;]=D:K(<<RFce]LSSg;[LKNOMgLB<VC<#N)J8BH
?:cFZ0I?0aa;8(IT6YEUV77>[O]G7MOQ&,;Ycf(G,-#66f-&>H_;4<(Q-c]4#7]9
+/A+M-W,H@gZF8e(W2BIeC&a]MNSD<[)Ua);\3\#-\MXbd4,JN-4)2B#b]&&NNSM
JY(#G?(+X__??<bFd_W<ASQ.f.[[&A[8)Ya:aE(cOacIAGAD18G/UN&47_Qb?95P
J^d6FaaUU:/KfVT0]FPM10J3eSFHFPYfLa-8(I33fHW1#?+<f/4GU<SKa3dcT_2>
CBP)2M\63VS@c/+Q;M8O0::;K4_ON(Rd-I=+M0A=M<3E--R9T>KPU-Q20P-8GM5C
O0[;R\G:,4\7U6?bSgX^<&RLO\R>g358GY?.0QPA_E](E+YM9VRB)RP0;Ha?Me5]
>gG[-GRZ(O_/C#S_V1,FB,2S0E71<,G=<_LS4C&SP<9-HDZ2Nac3[cDFIZe&^61#
F(VfBaF-6BET9P_+BSMS1E).MaW3S^GI]7J?U,-I<YJ@G:,:gc1QV^VUQJ5^[6MU
B@/YWT.I(5=-V\,d,MTf^FI<^c9d_AI66d4.(eab4:=^XB,S^):6J>)XQ>Ob/HQ=
H3=W)Q.=(-+&>R&E#a\#/RK_LJB1.?WP6HYTD?O9Ye1C0e@&b0:#T6LRH&XYE^ed
S/G1cY78<g2,JNL/PK^#1_gUUTBcO_^-+Q/36fP96[]+IfW?S^@<863#ag]IU,?d
?YTd>XC1\0M1O5D.XUT_REf_..NEWRF?O(K+VYFE\M_-.&0_W.@0gP5]/;1e1EN.
e9J-eN2S44(DagIY^Y#bN#5NYbU=^5Tfe\GUG>WARD-AJGBBXRA6CBaU7-0e+)d4
CA#3AcKZ^D#\HV>YbP-Y&=X6,Q296S@;1\C[c(ObW&@3G#<cJ7fNVNYCC3S^B5.A
DHK[;5,@e:)G3J[,:Z.QO-.Uab0E4]_V>?N6L8DM8PfXRc54P>+2)J\Z=#I&R-D5
01:^L[>.ePJ,V^Z3P#>B+)IQ/,:MV42D<Fa28,)d&B]9Ld94CR4bH0WVF_8-IfU)
S4=bKP\\#7a#HD=C6_E2[&(/3LYgOI[XB31PD>77;3^L[F[fSPAW8N3[GWAeKN@B
\DE[8,\UAbb#OZG-7WDGQ-eT/P@M54I:.P;BA?(0J;YPM5B0gF7F<Nb2)Of&D97C
MFeU_4#LG;W7eB-T5W#,H)ADS0/\Z5,b.3cP5+F/fdR3J(80f,4G#Z.5ZUTG?GE>
eNb.PUBXPK2U,-2.[VBH2Y,PGeG\JA+)7MF0\EAT\H;]D/8@MZf8c[X?Zb=5]QO^
W\A17d&#D<4[/Ba@8g9@6bVO9TMNFXO64c^a<)S)&<]?@5aG(\VW=>8WOOaL\;B.
=9.Y3Yg/7OL@3IfCS[KCbD7G(Z9a0<<@[UH8C?6>8+V+=)9_aP3Y.+cJP6N(=Nd?
8Z)\;@]=(B#d8NRc3@N^T@;]0<1cYNUUU(B]2GH\c/DF9#MUT;,Cd,HBa4ZH\\92
[Hf<0AEB+OM0>_3HX5J^;2#;\;[:H3f9^(Hc.ZBPH7:R)0Z&(OFGH#.)\+\BT7V1
T]34Nf(df,6f,&)Z>HW5DMcOUd:TH<ZDT2^S]3]:C,6b0bWC[D)V9=^0Vg^4aE+c
L,EOSc&g>7,R8YY[4Z8O:.fX>SHDYYM]7/AN/)\;P-g==8>)FaSZZVOSFYJTW7V:
[E+5:cEgUZ4HbcX9C]aU1g?_HG=fcB?=CdXR61IE;E-De470ZJ44Y0)g^64]TCcT
#47=gWUZ0#B]TYdV869NOD1L^(I^RE+\5D:E<]4L=Cec-HVDAIedMK:X<8N/&F<Y
6NRG,d+-W/BS06\^@JAS1]2P[FVSe=1f4(f)XPWVfKI(3]-8GA;&_6[?,_&I:@A8
(@9&I08-O/=&]cBfSC>WB9&Ed]<Rf_9-@Q6V67f3X??f/T.7EY(?IdQE-OCSQ.DA
dCE@bIU5EOBf/CA1L]Ec2M1TJI^WH9#D+5Mg]eLC>\&,:;&H0APWPf-DBBQ\-0g4
2X/](P=E_H0,<JBP23+c5AS>3RaS9/G:8Q>4]]>DK5@;DG:,<.TX7+[TS\V:]\1a
>g.HQ7g:/WfQEIGBb2&f0Q#7S]Z>7^2D?>D0P(J8e,F/)>]dOJe/NAF<9P)J8Y(L
SB+Zf&+/0@Dg\d+e5a1e8.e3:F8LQe)G0H1^XQHC7(d):S:/O;YHG9.ADD:EC#F+
G43J7@RXBB[ZD;0RVH-&FAgO+NPW&M^A[FN(JU\XP>Cdb?\W4P&Sb]52Qd;,LSZP
TY8\<JKeQR/_)65=&0_aMUOEbX_BRK5CEeY--[@Cce6gSAQVZ=6P,b:XE0+5B1&?
?ADHaEJ,F9E2HgB=X[aOZb^?,d8PQfB7^(BZ:+;]]B?/gX1L(=+;9U]DcQ)+d:&T
DU4bAP,4[[D1D6gLY#BaaY[JRa<[UedS3+(HB2WDB/B;d,L/a<ZA)MFcAR34Yb&8
Da@)6RfUK][=3:3:63XW6X[-&HRB9O8PI2CWZZKBGbe<4F=aDc+[1]/TH5:+gY/e
H2>JE\7WT(IU>QDUg2C;MYDU1J3>>GfZ//#e\Y2daP3.Qa(WRR8H_PDEJe/5M2G2
Of8LU>JW\8F3,eP/)],#FG^1/7)/Y]Y#@Ra<5bebaZU(JJDC+9YRSTE,/8G?:W\<
K\ZODb4\P2JK+VR-?e^J/6=FR25WbJZ=W]7D5&;G)K_C\&:d5_UWC452DN]2I/9/
F3K/S-Yd_0(2P8)HaSGP8\7.SdAcTPC3Q8f3OQ,>0JeJ._B]<:\:CM#MEXeJ@<.F
@8@2Kg30SKR[f;ITXd(=?g+dO47<2Z3VZ/6^HTX73ebNO?=Rf3)5;^cB845(R=7J
M1PdQ6:9.d.Q&6XafgcMDB8@9F3FOYS^Me[<0=<1=?=F7U\)fTcG^ODED)0,dO33
T:a#WbT/CCMZMSg+aQ,0/J:#cH^#-QONUQ:^7:eGK_?=N<Mc=>U<F_1PQKEG2V\,
<D3II.gZ79M(&2FJa_Zc-6R/((f,fXZNe<FF@QQ.YQVbH8G\&:FS(5ec(1f+X6=.
OKDf2ECfQ8@PECJL)4UR<_D..FfD>(6_M;?OWR8;(b-D06^@Y\Dg5/TSGZP]+2F?
,]PMb^NdQe@9&:]b+W9NAV+OTW;^,D_L7<TCdDdE9D3P)QAURUSEO(RfAXTWZPU#
K//f</UVI[F1K]0a15/;PUaXQYGdeV+cC82]Gb&dRBE67/<V(LK0^1ZQ\ga,e<^R
L<(XJM3#J3.Z/QOSK_FNE:1L(PFEQ1;aHV(:F1&LMO9NF#=ECC-@Y_LB<N]?R-)0
GT>a&WB.DK^bf8H6S5bcS@V0[f@eT)?g8eC#^[aQgL6OIMQMKXYS1R4YZ.G1U<;A
5__DI^O5.#BWVU1&8(KK+XSO+B\Nc)SPSG2B_Y;>,SNZRNd(>SD0T=GL0V6faL>S
-S1Eb(=H-PTD1ceLHMXE54UP#U5_ARb70.9)IMaB[,B\FVO#a)2(5;<&GdOLFEEc
E;^O?5)MZP-QO>3897QT[caAS?,-P^FG3e5aAa3Z@M#KE[9@?_L?MbA,g])@7R;I
#JDBT+#RPH+gZDARAM8NABW]Rf[cJa#+KB9(MBb\?)WZcK3COIKD>H[O.LbKVRd,
_^NQC-0NJ9&#gJ<M?\IDX/BD+@:T\=4d3PO+-:ZD?L<C-aS;,@;U?\]dPII,C)9=
dWDS-Sd^bA)P@2a_6[#W.\TW=_[ED<W9EZGI]NYOE_L(TeL/IYO&21Q#O=]Z4WYF
,,FMZ&YaU7f(?bX6-E.Z9:O8;UT]Qb_Q/T<<&J@853,N59ZNQ,3#S^0WgI]3>SOf
g>]EDWVfW+ZBI5B.;/DACJP6#QN.aRKNE+d:)06R]8=[&(EX:.4LHN+>10O&?2f7
GJ\bYW:#&ZL0FaO0C.[ZB1S+d8AIHe[IYN7;]WSI+#ba[(#QMD;>B\1N;Y[Q[D.5
e1#+=D^e2=@QYDGL?+d,HQ21L0<P5IM\_B2VCE#416>>TEgQ/KG/UXbBZg@9<_Lg
EW@GF8H=PeCPUA5bYM[g(J>M.B/08?_HDN5HL70?0-d4W=eQVb3-;A]Z-c4&-Jf[
&?AL6#P8=FHZ5)O]S)O];&P,DKPd^(=B7S<J&AbA?NQ\/CT\9R9[U9]8d0/PN]IS
K]41cefU(&gQ_FUSYZYB[;aO8d-8S<-bL>bM=\9L#G/7cKOI#B5SGgDf<2QKWFBQ
^WfE:6&3AWP/=H7ec>I3&#N:e2gD^<5H4&d\6Y-+IJ4cF@cB@<NO\E]5+5@S76#@
Fa+<WKW424S>39-V]:dO0Jf<_8=F3AV&?O&4gL:GTGg7L4<?O[(+AS,+:dTU>>-6
)ENc-<[#LWcf]T4Mc#QJCHKbRJ02/?f[S0bLS(432X<H]X_aFa6.XbgM4:T0a?eC
DK(LN0b/RQ]Ka34K>@Z3<<:c3.2a0GbSJZA^bMNK(.Uf52HE#dK2\Tc<#ab&J5Q_
B[&QM\6BSB.Fa3AFeW?=cD^aNC:_H)VO<(e9J:WO_DT?fUX#H-,@P>C01K.=N5d)
3OH6EQPJDQKZ[^?A25fB]0.JI:,N-aDJVcM.<f7-O;:(7@@KT.D/gA5BGYC0fWI?
K3Z[1aB<J@@gg?IM)(IM.WTa?[VLAgV6TNH:fNU>3).(9-?B&Xge<Z@e.A5b6fOK
&N/d?0>dJ\=Vf</;&W05]N.4\bQ3_SD82WAPX+:HaJU9@133V0dSaVG3f^>(WM.P
,2&8JDN93cM\6K67.H\WVe3BXQ1aB+EJS9TRF(=)0],3?1\PI(O;ZDFU3O9#dSI?
OVGQb[Lb@_+VJ&#a@S:>^95#7;OIeWWddCZJEe:bXPA&B,-MSEa\V=b4]O_F)\]M
S([(:>\BEV:RRA6RPd,&LV9I7FDB6M5.gIR&9P\b?1JOUY39^+?D5JeKR6MR;\NZ
\,>c3TfEB,J4..8B2N72#DXa0AePK_[,[Uc&AgFM4-1_5dd7K4<:>Z8-B;@a:P.K
V[91.Z4B3Ng5@BX-SS7(AJX;0e\4NKE?g3?TV?\J@=NKCGeL4fdLfe3\)@C<Wa>P
<e[]M4QS2aGT1B]6)4bUEGSC?Ag1NDgC13V,KV:1J5-Z\R\\dKF6a\.]TOS+8LgN
_)V@\5O2@0ZU\<c7b3X^+-8EVF-+aBCO&QGg5AH:D++6M)JNHWTUA/=[&71cCD^+
+,ZV84F/U-HEg3C[,CW_IO?#<361+^M@QQ;)(5EE,W0)C4\WVZcaTHE2.::3AAfb
:G45Q[@X,Wg;cY)>^ZBARc+[9B+=ILIaBL7Bd5O#M-+.cCH9b@f8&IN:ZQM/23gD
MV(D3TdcN3D5<.+Z>4P#M3fBQ5FOI8BH>0W4+:0\J53\XbEV;LA,3-KcgND1ZeW[
R+TLUJUIVYLS(3[W-G,V#@9RA.7]QC^Y42T_,X]=X\WO#a.4NXSYB;#1D_0,4XW:
^=+fEd,4bJBWK/IVeYB)MC:1-Q\ATT)EVL44K1PT3fF8;1MR3e87K<W.XH-d,82b
=9\c,S9WAQK#IWGS),f:99Q0eZ=d0C;QD/3^/7;I4K4?c^OBYNJJXP]=)K_RE(dI
6,^:RSHR9Ng(V/MW9A>9(:BF/_,8IOI?<,7,VegaD1^/LM&_1G:g3HJC&E.g>c99
2+3JEF0]T]@U9YGf:5:(3(I1<M[+5M+P)+GL+-(E=3[UJ8;Kb7TY4JF;ERP,d/C9
X^Ac>,3URFJTCWNeCA\(LV9I3&?_/^&A6@YP\E,d<OK9\NY=QCOH/5=g>S7TfZI9
ffYX6X?OQX_:)(9SHNPdFedEK]cUGCQ^HO;ge+XcdB(FM[0\-Aa<+Cae,..H_1/R
.@ddP1;V/F-<-D3,;T<NfOb,cCC1T;20E3W1.;):0M?cG#:#84XYAT@gE6W4LO<E
Z]ED8;S66fXBSIKV?BYJFX2P9d)/W9BaT[4GL0e7;7QEY<DZ+cTYIBAE,FA/>21@
6KLQEJZ2Jc+>-IQ6QM/gI@W9RAd-^(-&B?J.8>V(7B;>\bNBI&_-SOSH;LZ)JP9G
<Ab0@&=&#5E:+,NAQGb-<=/^L@^\&U.ZH&\9=/2E4.P+>/J,<;9e_(K493(bEIT?
/G^E,GUYD^X:GLMJeC@Y&G,PGCb_,>6dM]\SH8]J2Z=bYeFQbcKOX1(eAG]7?:_M
_TDa-D:A6Td9;[E>cLZX^Yf1F43VObC-F-7+&U6E^?0--026,^eKPBDCU8[KKfJ9
-DC9:W@\3eK.>RV4)[GB^cUb/-EMQa2B)?-DcTS_I](a9+)K^99NNeMB7P4YTUL8
1+Q+T<P73d76b=6U8_PC>3[JTb4I?4ZfHca>)#1E^9T&[YV9f,OWg1CJ<2dQ.8W.
,2+K<MK=>E>JE8>=C8U-/<<>FY1bRVH+-@D9Zd(WB\:4W.HPRS)A6SZ\)3/I9.7Y
JSK]QP\cSZAW?1D0(W82X,<gVaLbHKa2Pg6^S;QBEA[LcU6&GQX.T&5GaAZBV(/b
A[e(-R3#&((249KU7L/R75e;3a0;@AJYQ2C?1;Q^LFY^=:GK+@OS3[_=@GIA>4OY
bI&O&PZ#a^#_Vf4+9>OWM]+[O)]Z],WHTA^\57?c&IN>A.f_>/_d05T=a:e,)SMZ
+cU-d)e(NLKg]We5Q__-/EAe6g#]S::Kd,3&8->aJ>V?=gFO:?3<Z4#G93XD_;E1
&L&8LS.d;4e]_5K,eX+DG:>LYc^8[:+dFbNfE6(#?+]C]0@=f[T?;9\,Ue2T3(?]
):?YJO4T(^;,L7JVV[9GY4Q.Z=6XD:E+TeXd4VOTY^(,]Db8Wb;A.:g^]LgH#2?M
WLM5d/;;3R=;+dWG:5XRN5A,&D+3(Q2,2Ofg-4?2Z\+.)b3EB\B^;B^MD-L>C]83
E](+dE]N>.?]f/fb,Z?=9)QfS>\(9&eeMa;AC,N3:,NL^D][Z+L8:B:T>c&C02&5
Be_]gec\_?cM5YG\<P@;F:_5-BW3ZM]7F3<e]UNA-3,(>OP35[#&+VZ5P/)BJYS\
OUI0.L<?Sg-b,QHS0FUCUfV[?9g<.TfQX.](62)e7H)0?e_1OaA#dM5ANY99._3d
a4:S:;9)YCc^TV=O7G3,#XI?b>,#/6;4HOBeZIH>M6[_9+\-::C8#VZ5CFe+FM09
@]Va+K&.,FTT?cTcE6JaD45D-aD,W,;_8eHIf&V-bVD),cMXKCa9PMOWM4TL]JBM
1dV:+0?R6bWRDaYc<#a^B3KT3)#<BF[GP3Q.<VSQc8A+C,N3[\7=]V=Ce/4EgWKV
L,gN6LV</-8C;:N-b#H]R6=.QO@fV&bT?65;0TG.X3QW6U/F.06Lf#6KP;/c/G>S
8U/B7)&-_#6Yg[fDIL[1@(>S33H)E?HK.G[<;/]bTS^Mg<_S[X^Df1IaE-V&/Y^&
I.Zd.,R>OAJ,D)6OSMI?L58Q^^9<4Y,]HZ[3QeB]5?^RY5KU2A,P-HWVZdD<O?C,
FT20N8f6fFZF1[1>ae#/YbIf#-)29YNCbSaF6)ef)4TZbd_6F/W.9g4=Q7cOE#2S
^9FGL6,aMYZ4QK<F.,eCU2KPQC<8;^#-)-N6VKP&W)<^2V3-1/-YTJ6<Bd(Zec+c
+-(>E?48DTI1MO[Y<M#fATR:X6P[J]]O)(S6bH1/O(agU\J1@WUB)(DgQIXF;;WB
;:2a7O.0)6@gV9W4[3[R;_&a_[@DYU^.a#U/RC><Hb>WA0.Af<X?MEP/C<.NA/NO
G9\1Y]LLV0XLUT^UBEU8V@I_Z6a_4W5&c)CQOK;SGaFXcZNI-JM7GSB:^<VBCP<f
cS\QNDO_(eJF)S:@_>G@2AC.CCIfKOSK-,CJ#AQH5(-D&f)UTQANFfK#gC1e;+J_
a2D>[_=>Fd9FZ&</4+RXgMH]KG3FM_/LU/Ac41EMI_ac&K1G1P0(.9gZABBPY\)c
F>+-.EaB]9)E89H1(ZKYD<ZBWFYJ\M@dRHf.d?ZJFZY\51G,@D..8O\XR_49c0WF
4HX\FK1_EgB[g7;gQ]^0=3LI467UW^C68.WB+/9,8DYJXB&,Q]JM^V,bU95fd,Zc
DXN7JQ[&JFWf7,<4XK^(4g@X&6D&-:.V,Y90/g@ZN&-&=KSPGY1&-[aVKBd8IS]=
2)L><;IU6RJ4,E94)/Q:[7EJF,UW5N<88>POK,75_G):YRf3PM4U1bO8bICfUM&/
H@F+7a;cP?S)@L))][+]c52RV#DWMJ^O#>;-5?VEgTMf5aEQg/1e@/(IPAQM;e(P
+TNJO1]^S9Wb9B<XX[V3=L?#Y:#2GN-8H&=e+BS[/6[LX:)YD[b]bFEf]P@3Q[1]
#8?=-8(/:+HU(^F+<)X/2(:9OC?].Y6IB4)LQcF-V48U,7;))2C0SRTH:8RU;9A?
I+O/E(=X._F+GJ8CKXORb@/JIU;dc2aW;Q^N,N+R]V3-K_6gLO8A9ZCGZ0S=GaE/
?,Tc?Bgd33f6?9:Fc]aAGU<5FX.)-)5R9:P^VBbP\5AL)=,FS902g1)_8c&4J+fa
FP64;^35/.7G_>&DaTbadSJbUOK)BX&a9JFd@.UCa^gUI:VMK>&F1fS_&Acae5X(
/,ELb7AMZ6,&]0Q.FPG1D,7#?Wa/)8?P.92C:FOXVM;g7S)Qc&I\fL_@?-0K]+]b
S6cI-Vg1QCI?A[dfRE[/=HO#]^S<Ef7L<OfaF-e@)<389SVQ@G@AB>O7&60&5Z89
XA@8&^-43M5SE?N[OEF:<C,V2&@M3Ec6fX<T]DG>+@3X.RZ.9C]V07a2&\;A/^Mf
9c_V[8.L.0X:g0O9N[YaJV.d/]_)BHI).1E:DeM@/_BG.Z8C1@W\J6N0dN,L)SQa
=VVV12=O\RA2Y2\V<YMSMZ+=gg3XD(-(QH\H..-R5(27=b#MTIc>/Q))&fB#8LDH
NU[CL6-D\LS8Pd[O.I1II,;3g5,gJLEX,M)0ZN/UOEE/eY&7#KH]GLXL7T_S#X?Y
ca8P3A]TA26E)?K(Zaa3?Y)(b)/;0E9QF_f;1(K(Nf\60/.PHUa5KfG-O(T6BM9[
;8JD3W#[Zaa9E3K@CM(<fe2BO,LOX?JT@;.<T^9Y8gP?Y9L2=HXd#1.-SK#U@ZS=
1FMT]XO8cQJW/FTMOU.HL&W,-?GBdcB+#M50-g\VN^eGVd)ZV0e(]T/I#?,0T58)
NcP#Rf,93=c]9U:_eL+Z79UK\4L24=T,eIYJ?U>-&/RR?EG\+^T2#W9S5TAa]K5(
R=N(_:+XRB1)F-AcI=[Y+aXB/8PYKY1V&dJfPa:YE7X4F\4F2]52)/?Lf+KIbHbf
UKA)W,LPSaVg_E?PG-^^/8NMTRb4;ZYc(P53?QQN[<JP0ZRc;@/HRCS/KHI)d;\J
0;<>H])bRC&0C^LJ,6P/V@_TLU:KE3P->>)G7EO)D>6R6)7G+fg7=d_FLQa(XB02
R)E8Q1WX792?JeQI<3T+DX6Q:/4W+6IW-O8I#?d?^&:9E4VXNZ3\N4H2C]/[PT\H
TP1f(KN#gP\@B+FZSZNg,(g.bCJR3G](eY>KSZK(fYX4P^4T1>a;&b<,We]Z8g:Y
Q(7V9JS7fWUF)UJ4,\_.\H^XKeYA;ZWgJ>a_[W=)J#?KC]XSdSCeHZ\.5&ATg=</
+,,8gNLHH#.cd>:S+R\c6[AE:3/)48ZKe/VJaMIZRJH<F-8>/Q?&bF)H9_;;O&6=
R2#?7/&ZSCAV+<M2_]84^)A+P@;7c(Y:f3;DDJdf1T0aeU:V+XC>;7MbGA2=<I>6
N&&XWL:OM2^4F?@:+efZ@Y>537TT0:.K,2>aSL5YN3(a>,L6<Q8f85g@L3^;cgW(
-Qb;bZec2&N]YU3H)1/4eG0J&W2d@80R\.>La&9@3[27ABgWA.OTI&^aE=)J</OX
bTGg;?T=?/>=YYN88:Sg68TgU2ePKe6LZdBV?E(2?(S#(UK_S^Ta7VYI#KT9Y@VE
25,8N:UH;]QP&1P96G@O>[](W]TVY[bJU?-[B+B:,Q)1KN+_)M+OZX-59.1JG+#)
X-7W.7<AA&N\AXGTEPZSB4P//gZ7VMPQ=L-TCP3K-M-ag)VBO)8NRA?b6a/0DT;K
g:;b[QTXJN#)W:V7YAUWS3&P(3^3K8,Q4GIG5VBPDd6<;3:C]M9Cbg4X]0J4,@6F
,0Z94]L5_E]HACX06:G]2gJ:-+5H<AZ-^f>VZEC5MTUBB1KKdbK_NbYW+PQC)[CB
Cc_N?]M)ge(BHA\B0a>1/<3<PY9H836MMZfNN#YQI5<=X_MESeK:Vc_dd=D9>bf;
4)=)0;5eA.,6;9RddD8a9&d-T/bc((T^gd#1)fTBBKFU=:/V[C-R0FMGgFPfGC/A
A/F5a>TUbC3:4S.N8X(-KBb:HC((TR@-?G;PEO>)8^<X8EN(TN:;;G8=T@5,f0,^
<_OWQ@)P_cX,H&Q-ME>6_c#;(ZN;IX_K(/f3E/P_L+@=V;aN8O[I(cc&]I91d&-[
.G/gbY-RY@aW^2@@/ag,D\dYL.MTA1:NANWI>cFeG^V^CbRcW9W^<\3U]::VCI7O
]bbGT#C1UE:@.S(C^:b_@&+(WL(,afSI0\JP1Y0[dEgGP@#LY]48T/YT2Z2S[Ud7
&9X@+VV[f[aa2[1QP;)<cMUIH7[02[1M=WaWU3R7FcF3]8K:6MTcW>BPIF^UWR=d
=;CG--_@bO0[_G+cBD2J,eS&9+7Qf0NAMCa_XJTJP5+N;3+(^FR?3JUOGFPCTV5#
A6+)E48Q_GP.1;2;:+48?aLZ9eAWSFI5S^,QT-QeF#&e:d9e\?X^D;.T9VD(F=<R
4V4T#(F3R<RDY#S;S^3)-R)ZC3gAf(4:PgfM3S#0)_7BeUGgBPb3e_MTaYUdc98Q
H6D=aEY.<TF]9LGe[D6aN_JD8b0LI^Ug:H^?dT[fM9&H;W3YU?WVdQ&-LS-SNXH^
=ZS0P6CcA6J3EKC-:SI(Hg3[=;[D4Y,(QIDMV\bd)1J92:7(O3)d849N45W[CDO+
R6CKF8D(Z0V/,FZ]ZU>g9-O;5&QE-H:_PMM3]6@(+==dI2UbW.X;4cXbOf#2&-EX
a?B=HW=0]:H?,E4(H+6Ie;9eFQ2=GO<gHKC1cT+,&7Ye[_YZ)gN@&UASB0;UB,=C
FUZBUO#Q>0&K-WFRR>O_3,_@.,>@UED):XA(b?dXJe=N+aUPN.:#X,bD(I(P^5CB
:Ea[9#:TR(XWCeH/>6fH16D3Ee(bGY^.=S_&/BX.[-cbG.@H[7\45#<BeJA:QVd/
38=gMf>N\X+UW=)Wd1eEHEFL.d\^SMN=(62TE<_ge;B#K.W[]5a&Pd3Bc8.9Tf]b
B^L>0DW_G&bX3g?M0>RIP9-IR)+84Ka>)BCX0Ha3fYcY5Od[L@1Z#.;4gU8X3>gJ
C:6.L(g@-2F#G-U-Z/208b0.>W(.GM>dJV=J;b0RU^Y+,8dV_RMTb_g=NI5)PRZ?
\NbMgbHOK0VUOMFbY3BcD.,D0f0PG@-5GR15cU]f]9^,N@Z5LW7AD3QgRIVSS)\K
Q#/83e9Uc]_?\fFgWLg<dM<A0.;T_ELgSI8VO>E.SLL_d0b@N>6dVZK->0^aROUJ
2]\>]EV#Jg?Q9WaIM-8I7?;@F(=^TK0_Wb<:+8fSR2bM=LJN7G98=dK=SSM1IcKP
5Wd6b)I^&:b5NX(T@Vbg/[;&TXU;1f\@g&&G-C6VLcE[f2QJ>+;Mac_R.81F]6O5
+-41WXF\L<_F7f37(3JR\B_;W-V+4DB)A5#,]>BfWbfB>(+W^a;7eU(N)W6=U1<A
YUS5@S;#;>S7RIQH6:0JLIS:IS;7=Z1.[M]Ee>24P@#L2:[ITDGP>bK\UOUVSPQ,
=V-EPJASdUX;@6]7HW(4M(0MHFc,Z<QPT.e?[[fEUEJ?,8I9K3O]P14=)K,4;EY(
dX9fKMfZ=X]&MdILXC/^DII?YQ-af]gbIHgK6JgY0R/SG^ZT.:+69(W/QFJ-?I45
DbZ=;3KAN6709/82/1\G2L7N/YP-9Rdf(W36AaRe98G7F<&H?>8-UEg,MLCN5//M
=,G2e-M-J^@WHBUWO>.A3C1BaG#@W?6]edEB@?US1?W7>FIBGUK,5J(:=LCc^GRK
L.B1C=G/+,(2KOPA\@J.F:bP^5&M?[W10<BP7C03&QeG,9L>dcX3S39/BHFVWW@6
fdBFLgF6(d0M3&/d^aKLR?+F-VQg#+Q7WU^e604>DE0F4SaB\>M3]U,PL6STW8@#
8b^J6LHTf<WAY\b5K)9R9>FI4=/[=F+2VS4cQO]QK56#Y.OH3/@^gL0)-[f9^SgW
ZBCd2?277-<ASb6_NVafDEO[Aa,C4#RTZ[<9YN_8gGedZd6W1TKPO#]1)LeASXR8
O->QU==c&L8K1-971+01.=F9HTY35V>1S9,Z46NAB5>(5ZgEK\[YX^@Kd_a[R@L+
>S/UT&ZN5Tg#&6P+A[W90Z5KS43E-KK_EKbL^;+:AEO?bN(=\.CP3W)O<5NR[g.H
&C0@g<eS45BXHQ[+3)JT9Y0IJc,F4aSY0&VK>Z(<U&>fb==2L)gH5a&Y#^G]FBN+
>>K]Z(BE9,Q:DCY33-d&>?-N)KO4Q@;?P?#<1YFAdHGWNVJ[ZSf.S28)3QfP^ac2
FB&JgFELaGaIM&\N?5dB^UW/c:8#b4+=a.9,DI727;ASJS88K1.L(U^KNR8#3Q9F
RfFX\?SBdM^ZgX5U]#2d^R8#H6cT&P7IN+#PbY\B[a[I[]UYX1LB;DBSa8H=<D3^
1CP?&d7E4L[-,aV42=aPAd.bU]d_5U]gWcMga5KQe^3efUXW@dW)H9=(b=8CJ.A-
[EKJ1UK7J@^92_1>6U=:A7ZN#H@;DI+)G^a<&dXL+ULDWH)J\)9Z-bSOP:].b5[K
Q2B;2+7-6/Ya0M?5<P@[>ZPV1B;9#,0@N+[^G,14</YNUX6SSg]^9D::VKXH@Bea
IT):,28+G(-,PHIYV33M8LN>V_Y[3XQ:a;Z__R3^]bbC_c4bDWGV6g]NJ33=)6G7
/U0(IM16(g:8/gb_e,^EbbWJ8TQ>VU=Q&cG^F(#N-O[-OW1B2P<-5>_LNLC\1=<J
a@CG2IYg[eQfgH3fRA1ZW)<[H1,K]3[f(^I_;cZ1Y&6GU_BGgP1&NGUMNe5aO=18
U/&S,(BbOaQ&PBdc+1Ka/,4X>37.)ZbS[RQH>KMT,?:/Y90f?15M=UYg#.1\]6ME
O7b6=Z3;7:=-DV,:5QL=^IUU?>VYM239K]IdYRZZ(=a]7Pd<KH)@MKHN8Q:\9&A.
6YZCdS9D&.>d(8?<eb_1A+AOXM.X146\C-61a<Ac)e+IDB=(Q+e>PgdQW?C?C5O&
5Q-JXG+83<9WfO^,&J#T8/X:Q@A4@,E<W)8M9/+80JY[b008cBZY7-UZW4<EU^C_
X>W=QG&f:QR30YF4Y3Q_[8U#4;1?+(a:K<K/;?gM[JD=J\VE+:;RDO+CHD7R6dIX
.;SEUA3U1\8Wd+E@6&7JXd-,4G]<QG^dK,.;JKE2@[D<NUaaV>[(?USa-+MCRW=X
KJB[B4;X#UTf-9g])/&YUOC[([PD.&+6aRE4XZGZJWWIO9=;=e(>MJ3/]OOFJAa+
,C#\+[M>AP&WXX4ZKAQK#B>;WO8f)=(7,7FT:=K8U[ab5fb-[#U_C1^3#X]]OT91
KaZ83MARZLBFJPaF[UI,)Ja90K[E9)QFOU&EXKWYWLVa;K_&5P_23>gE0bWC99[3
.b<CHOTD-FW_FYRcYE_NQCP,+)OWIL,G>JQ72aC7ISK^J45@5#<?LC?#@N^(9KLV
=A_Ha9:60=;4dV4d\^J^EZ@cQ2dB\M^+,A_QT2bL?.b?^/a)^RZTaXd+P5FB>c8X
MMbcRW#aV88T4c01WDZ=ULC@+J_5bdDRMGbN&J(#VB]DV7@>+eI@e8QQ<06M^(^@
-geN3QD0=Z42Q4:HY&;5e)=>\:I3cDD\A[\==T_G/=O@NBS?^3_e7NEVS,AH2TU/
#N0U7L.cR\NPTLPAMgW@J\_=YX<+]I0124f.df<,:\Q?_5V#GW=1ANINQBB(aLY_
IB@+]d);fdWg0e2U#_R#9@PCJ7^e?[2H+dfQW]+dcKTa+.9NO\7+O>G3>J=8f(RT
ZLQ7WW37A1BECI6O94/NHP:(e]PPX9OABNU>L1<RBTG>6aEZ5#?V3UM4\5YP^]_+
&SM[];JSc36_(e@B#D/9VZHWYK0Y9TEF-^+02Z9R@66^dWP(B92gCddWC\B3XWH>
D;QXAJ,WV<^dbKV7U3\Y.gPY2.QG^.Cd<V1PT9539d:gCbXHXYcfYBKC&#a8\FaJ
>^H;X5K.5d6H^);+;?C:baCH@CH?TYEHHIFI?E\c,_NM/E5GQe3_3#SJ.f#28Ee\
\Z@@0^>;5(<(LbgDQS]G=2>2I(W9Tg?Q=1,J@@dc=Y(+JOb?Dg?Ye.63QZ=B@UPV
a7d0;_O?Oc/MW1HdWg/N+JR&0+].>TPd5&fS23G[AHRGB9Of#CL5YN35b3e29dWK
?;W\3@;g6GTTLXR\e>7.+3D9?#>24OVBZ\=PgJ-@OCaGb=b5L4+E,^=f&cT=>M>M
XPJIU/9];WdH/?P^B(-JEOTd^gYY/7;13O+[fAHfBHD\c:AW#dXM&beB)DQM(AZ<
JWag@a:USK[I1W]\MFB),0B](:.YXb=G;E9^7(e\SF43RS,3R#?^.U.+f3^<X_Mg
+b6\_ZRE.J@P4&C,#g3]XK+/QTNQ4@?(4ObV.+8c7?B6C#Y7?Y>6F.UJ;UcK]3W>
O0bJJ<@53C,(GLZf1.Me3GAF&,^dAYH_EQ=E.G05aO<4?a-FTOXeOEY/geS?S,_J
9@0T2C5Y&:8JQNXZ+WLaf(bbcXB>NKFZ28D#=;:_=]<=H^DM0dA@eP7XLV=;e9VW
AEgDf57\=JWVcG^:I.:.Wc_#N)79-FT=aS=Oea:YB2WW>SEOBDV](.CdCBF]<EI_
>U4)-@We\VdEg15(NHHHPL9.4\7Xecg/f]I)cT2VNDRY_)U3@4.WU&eG2_4WebL4
OV3VK0:[8Z_PGK:-a.A@;FVKP,G;L((RPP7XPg[K[L\]-JY<?M#3K[0S1Pg@X#9b
&c--0QdS:\(Y^_b/_4F[CB5LUN<5<T+;_EV^(C@Vb8?gD,WB-2?+B_-45B;=H\\]
K^b.O?0@g2H-G)5EK0SY7:?aed^g=M@3(ggN]]TA^\f[275Af/-ESAU=FD<cM?[<
MA=1,fE8Od;SQad27)2I@I^9DDQ<LD6TS?AK/eE+WD9L;=gg@Wfa0>A#GL3GUB_6
2SHXU8ReA?9)Vb?0IP@1(PO.)d1UdAEga>:,c?D)MfOdUN9<e6+3I-XcBY;KBeaD
HRE+F1NG@>W26_NLGV1:S?aT,;B&L(B.6-E,-&Ff0ef^9??g8>4?VVR(0A/+SY=_
G:,^V?gLX57=<O=OLHO@W^dNG.O<^.<7c]G)V>G;Z&ba7E<6?HJ5=WXHDF5cP-.W
@a_2[)Vcc^>_NU9_SbE3#EEGSFC__aEY\V_Q(IGRAE(6(2BKU5OH4/:@bZ[-bfFH
Pc?5OHC5,4KcEKL]S(P.=:Q^4?MgTf&/BUT9aC\Y0.NQ?3/g<59dG)TbA;]Sa)\@
0<6]Yg5LMF@#O7N39\DHgJ^gS>H&2Y,CM^e_We[c2^=APA<B1+?,:O,]b(T,)e0;
ZCfHFIH1\Q)Q0^]Y+.Z_EIG&M@Y1-;A[AQg6a?6JHB^4J=BE0T]0IdE2M4GE8>\Y
/WS[0XFL_/He\\JTI@^e3/XP=?NA,XVY;9G;?X-SeQ>;MSdLAD&Jf0F)5aZ7WH(/
F:H417JY94RMMc9I=;O7].];;A\)_0R:R,QN>Fa#a2P8M#2dI0N:)LAV>d5:]-5B
<:T_2#+E2P<7M^f/EV[567ZD0^KN9?;Ze^_f<[CaEH?NKMOW),#1SS-e\0dB62/f
/;Z#dR]ebYP(1[FR5Z83UQ<FR)-8Qe;BW:@R\YU2bV3]3Ma?<51BIJQ-^OSO/P84
\&GJVa\<VNS;)\b:U/IBSS<X8+_IPBTHM[RIb4?=cV9MILO_+P@FAXY6#\Ke&K+a
F4aGAEgSA.ODfK0W=3Y+1VJ:<4Mg,M;<8T\&B1U(.fE+3^.^OB#RW9SW?.a#O\,F
TU41_#MEK4U=RB7\1VFTRd8.&JH/R1H-2W(f;\:S93a(TY^L(9S;BQ<F\J9D71]9
D1_1^cMea2F376c+&9OOT(;^V<&d5,RT(dC&O\60O_<;VO?0P3NEDTd(]_MffAU_
:,6cbEdT1bSIBE&(&1AB@dWCXDRW?Z6?cVC0P)(E+R#PB^3K?@2G22e.&M1dU-fO
?>5Q^;3&#JEK>=2GJ:J/.Gcd;Y\bL]?,.IUe-1//fD,dFEM:K18IF@d;20f#8(^a
-4MJfEbO+bd>82DPKKDK8Y_D9KIEf3^68Z-/O#WS&=4T+L[9.eCW_#(daG@^TI,E
>@P\9RJF:.)(M-55C/P;Z)M/ScL9[=@:BYI80#<_)8eZeP846]ANXD?fdL[Z0<Z[
(2[b6W0-a6a&W(QaUTaV28Ig)F(8BQH(U>TN2g?OXZ&B(+.8KS;B,Le+Jd5Qf>ZZ
d+bA)UW75Q-0&;bBZ([+=.;)(\KZ@c-2c8<1:7;FE.3/EEE)<\^#_:)A:R]?&Rb=
9H5@Q::OTL_Y9&@I+597@(?-ETDIc;g#8^(J72a0d:=)?4=Ig/4)H:aDcTA&+#4a
[LRN[HJXH?Z2B4=1KV3@34af/=bHH1FgScV4]E0DWf_>J3eX1VIVD>46K+Z@Vd3N
P8g4=9H[R=M80YXA;;Z1+ee#.N1_3baaR:aR[?a3Y,1RQ.BNK:Q_HL_#3]6T+1.)
&FABBb8RAN,U53-Z5=E>SM[WY&RV=[MSX:^KDUQZN,T(-O0=[2^19]:BV]Uf?f/:
XLSTX[Af]+[5JIA;^V,H1;<-<TQR#@FBG5,71P\eC1,78?2V\a,f51+48DU#eN@X
c)R]e;(SRQ^P93([32Q2a5d:R?dO&9HeVJD@BMGTE)H9UPX1,N9fTWX=f&?^E5T_
U_>U_[?bM+TBcc#IZDWKSQ<#fgg0[C#V0-1<7D-99(NNPQ2WCOSCf_G=Kb]LX[AB
DFd-DDCT4JV4N4S]5^Cf;XL(bQLI?ZgTaO66@C1bL#2g<.]V@U-RDE&)(8YPD\2O
T^fOa:&NAQ@DCK2_9>8W\>7f+^9F)cc?7,)KA,+0Ade[^AKVB?+((Y8X>d1DaH6,
H@-MDc]fPEJG91\SS[aI#/ZW.6.<5HWKD&KE2bYeO=d9R2)AI;bGE;8ggec_8=eQ
9XO,:fO[>bf6G/4N-JQ0Vde6&A]UKR\aDD6S#@6P,WcCWEceE;O37;S8O^^A2Bf^
?<P+==Z;Ra:;;7AF9c3-1\(-1>;EH1LdXTf6#?F<ZGARRB8#M3F4DE&[UUODS+X0
I0fIUaLVZJ&.c&.SK(70@+=A:3)BGc&.UD9G-YUDX^TR6PaC+UDf&)T.E=_T=G,f
0;CLG+KKKRKWB58SGaM\fI7U^LFWN]5RdZ/:WC<f-QX<:@_Y(1B5&7-Z5REOLVJW
-A/V0a(6UNgc_<BQ43[HWQYe52&C(-^[^#@YK,MIX4<4B&A)6.U<D<SE_-A#=?V<
I,?Ke)TRY=7(CMDfBV,ZeB_6MW;<4Z,Cc&+(,gJ4\(6c^?0@2;53#2G/@.HOc/8+
g60M(G?18O(?O5aF.GAL[7/)6QI@/c1C.HWG35a^aeV_<[X7J2T4/fHWJ6DPXbGK
,4RT\/79MX?@JRY9YXT4&C;W8VC1^I6F:RNP?Z1&BcS,>GFG.:@((>YI+3#)TTN>
SJ/G2I5UC0b?((0f97\)R;R.XL4..5/f25(8cY<UAcefEf/@DddQVC_aU7fJf&1T
:6+828ZRaWY?XA,9AfcD=,FW]\_;.Y5&.C3104\a&Q8<Y^,,V38BT6O;G-3XIFK3
=&CH?F?^G.>O(Bg/g.6aV2RY57#3VG#[)2XHVP+4g)5LX2YO2,,VDDfX1>MQE97X
01R<4OZ3CJ1=.OX(_F<XYZ<JNe7(6)@]gW9H)558DXI:R7I8[Z5cabA#JTMX8Y2a
ZRC2K=@376XT6?5Q,O4J)O<J3$
`endprotected
endmodule






















