`include "Usertype_BEV.sv"

program automatic PATTERN_BEV(input clk, INF.PATTERN_BEV inf);
import usertype::*;

endprogram