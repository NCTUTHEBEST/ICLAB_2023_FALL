`define CYCLE_TIME 10 //cycle
`define PAT_NUM 1000

module PATTERN(
    //Input Port
    clk,
    rst_n,
	in_valid,
	data,

    //Output Port
    out_valid,
	result
);



`protected
b:D_@3\4.U^cKWgBNd>T)E@S57L)Rf:[[TReB[@:RObO+;+D]cH4-)TMJ_PcEK+:
BGXPR9eCPbBNa-d<MRe/e<f=<_3&9#L^?$
`endprotected
output reg   clk, rst_n, in_valid;
output reg   [3:0]   data;


`protected
>NU9AE3X]23Z6gV2c8>=I8.VJfORXL+?B1aeH+E)c=ZOX]E&:;^;7)_4g90IWN@N
XWQ:^+bI^7gDC2A_=-6GDP+]@WSg=<\-/[S_#L-&CFGOA$
`endprotected
input         out_valid;
input         result;


`protected
H=44aLNgUUX27:.MK:D7[KO/d-c)OK&#aV;(Z7b?2^5&4U>aL^E>,)XZcf)4_6MZ
?9CEb>,NA,N&Od9\GR0Tda0J0W=9d&XO\O/]H#L;OIL-Ha#36XE(_aP+_eBZT39#
WDHMPZXT85Ob?_GCU/@CXb-L#/I+;&U1dcRI[KH)&6EGJLW_([43E/IQdccJ1<[<
=7C;.YM9A3>JX02XCI(MCS?RTd/MY?SNgK3SRK.#QS=EeAg-ZPHI)YF8&,DeURL:
[M\>.J0[R&.Y=6S=41W@-5aJ]O8Y&\FWfV&EGGK@S755?]W_Wbbb/I>;YdS3/@S^
5ZID8-@F,Peb,5MEBJ7]NP(U@8/S,?MaZe+;@D)Gb^Z+O05Fd0G>)7LbN04d[=:a
R.b4;))-\cIcA2AgA[WB2B20G5#4.]^WWS0Tb(_MKgT&Y,D:((VOP873QUX-;HS>
74?GSY8GKWLf7-)/Bf/VfAG7?.N27ab#R>/5VeQ@-::PE\EB&=NdWC_E-UOQ]RT7
CC85L8EWIaTO\_3OYCD4+GdaJGTSW1:?JNbbJ.B;\09KI<?\+&CK(X)#I>44KSe3
65eA]MFHVM78\=8M(cNcf[D+ce@,765_-W86(2&4Q6@/cgWZGDLW\_.Z)Qa4([bJ
[Y[]c,L.GEe^](?EPeWDIES\YN1I02?g.Se;(SUZKI;.O@]<E>BR5-e)\_H^\#DK
XVN4]LFU08d,C()9Q/@LE/fULR8[fe:d/,3Q35.^25E^eQ#N)A/I0(gCTd1WE<eL
5eY17P(;6DH&gN]>Q7F?G9OUNO?&6@ZMBO]?Z=3]@QTX.BX<2H):J1=fY+_4?&Cd
A7M62B;7R_VV5O-PaGOTg-TZ\S1)aRXGW6fH:2@eBd?17dR@/5fN9AAc1JPN<G+[
OZgX9aM+YbG)B\?0?157]F/E.D;_8gV_g;eQD#/PO&WN]1FF.0Q:R&Q2/(D)<GXP
<aTB<cRPQ:]VEc>R0LM0dNE4RA/U/Sf?Md6d0?W65Yc8JN:Y,/4IKTSZP^=-(++A
8R6F:>5&[dIUT9[Z,a#.G2(:ZQCGWYXdgP4V^G7V0)gB2:)_ULNbLDg4_+?U.68=
d0d,_KNE^SdF&4-@N5TVQ#_(S&9gBf;]N>e#OO5.(.\N:<AOSA.3^8dgB[&YVd.P
SecX&O#@7e:f-J;O:8WJCg-V,2E^21T9M-.WG?P-@9A6g<0_35<NX#R\TW#QdEa4
4DS9#Q[.R\RH6Y]?6031bM<.ICbUWN(GIC\BV[O(@MT,cW.9_IL>./P7@/2=K<Od
M(BEUe_B;5^;W4e:T[6#K8<K[J1bOZ77A1.?19[QD/+)&/9Jb,[.dW(#IM,;[Q.3
ZPeWER^)b9g.]U/=H4C7J;=+(6Mc/6S^2,JZF&:c=@e1D_/bC7OO;OKT4bAGgbgO
RF2XWW+X9</DE+85LCfC)fZg?gf2?eT\ENeCbAYA^)U77IGRFM_gO<[JVOf@D[VW
&XVNT^)L#d7,=bB0#0ef-d]JcA)4:G_?N>5TOeM+RJL<[975WF(8ROS)V^ZQ>(ed
0?^Ue:Ag;W<I&3^3X9?O-e-b&@)F7S8;;M<Y0c)T#Te\9cWX6GJD;L?6;bS9+??E
?WCF2J@B-\5FJ\_>49(AXcBg.,c1OUZ7I?2FcD5b13M\WQ>M,X8Y8VT^&[X&8eR6
d(FgefB6W72Ja0M-bBJKIQEf/:,28QfYd_3\+DBMDg(3QJB,Z;#]:,2M3[=B=\#(
XI;^0B-&UY1K7+47C+=G,WQac-4f2SLdc-2JcXCg=S?;X=IKg)Ua9d#K^0;K7b[@
IO]?D]0)C1&M4QRH7+/c1O_VeO<[1J/.1NX)M8dd?@(?TY=K,aL^A/\/2e9FDS[K
CU;E.XUTe(53HFfc24M?<C92ET-eZ?V.V^X1c\gV++@0;1ON9I-4g(e.FJf^YB(G
7b?0fcD^3:LHMPP-UXYP74-RGd@bME@>3(b34&^^H/BW3cJ[Jg25,F3)\fU[Z45\
ZL72016[/2Q.9C+NE7ITBL)?C]YLW891[,3VOZKc&#f1@[1+9V7b(TN)2NY@bX6f
KYb9PW+X-;O5=NR+AT>[fZd;7U7C_;Y]5/-V)PH[ACTU5:PfXK:3>(>0ZXB9&&XH
+4==.QDAOAHQ/RNRe-VY^GTEM7]Bg5EbG,X2PO6)^AVE;9Tec/8RI>I8KXU47:&E
@/G7SUTPQ)OF.FKD5LXAU@WA>9EOI&MD>IKQaf6+YEb5P_H7d6bd90E.<3cV3]:I
PcN\QA>^M@=9]EE=\TdPAI6d>)V[V>OVaH7^@aSZ;Z\>0a>UF,OPKg;<LD_FOYCW
aOSYI#&&[01e/SJcAX&ReNf2G\fd-ReReM8EdA-\[6:(:@g>,ZJQg7?(g]Y)(E[f
d<&+5?&]ecXN30[6IPd/-H0TI&54R:(B9@IaD)f@+\OB;_+INBU<QX>ZKEPN5Ea]
aW+d:O6#VB7<E>G]WR1\1++VA,WD;S8]R&&6ZG<;_8EM@7L4Nd?<\N[TE#Z3P-3K
[NQ)c/1g7e;FFM(I9F\5H73,O-e^0/NP\3f[7R9T>&3/e-N\\CGF/gVVW@LL?A(P
:WH@TT9\(Q,7S1ZPMGS<dJ2Xe)63PKLbBe6ZCQ>5I_PdMSe?a]X5PQ)dg#T-(/?O
MTe-M?X??F(SQX_HS&Z2&a1IFOZA-=d81.Q(]JD6Uf06YKZ;K/@V-VK3d,R&.Y#?
]J&@TTJQ-,[f7MJGC)=-@c0VTYWgG50-3X:/PW(J;dYR;RL3_:&a3OPT@NXV0R>>
^,=L#2b:1L-D0X1&aDI5R:67.0Ob4<9E>UF;MR7#6R3=X_:2FdB=B.7Q>e.NN9bb
]G4X1c##5,+=+-3CW.<(48QK-B(KdWQ<,7<N-3@X=).Y5A/6,4eeMOYe6-Z_SaV_
gOLZR3.\9=B7f&3=O[fOZ[Pc:#GBJ?bA8,(_gZ48SH0./91aZ,F;E@KTRd]Ve&eH
4T&IM\H9J0^&(B,gPg.?M6Hf\f#2D^52-LV?<C;\<D3bU<8-(]6aLV[2+9(W]L\^
S[N9D5^&[:&.?V4aZL>H?+9JCS=a7FR_<ZL56KE^E/AIZZ3GPH[ZN#QA,;9#MTBg
IB<:ZgRc_.:V@_HC<V7V&Ud\Kd-9>M<6;^T0=/aSN2KA8)f[>JAHZJC;eF_D^RVR
LY^25Ha(2ZPQJBd6Ud=1a6E80=R1J-X35@R.-76(Y3@BJHA=F1O05<9@F(N^@3Q4
:8:M@N^.N,C_TG]NEK?W9ITMaJ^B2M>-O7Q<7aeU7eY/QRXd-]V2gaZ1L/:g,K&H
#U[&[T@>T+/\&f>PAVF9VIMR?JHaM[aMaM4Y0AfUUb=0\)O5@L^+8aOQT090M?1f
AU^MS2>Q9feb4>:GdfG=W<:b>6BC4)K(2UPR8U7Z#](b3bF.2?5TbU,-887=F3Qf
Y8H([FBQbGON7[?U&P)XH)<E@?YSN=+;42^RO:0^NDC#NW]T6472^aPN(S>C8b87
VENT,EA3H1JPd;_R59c2XgK.SG//PMdU@Ta0AL7A)Y8J,WaDgDcQ/dX+38J0aOL0
X1_)#,.McLS8NQFRK?40;C+,UAfW3@:I_6Rc1PIR8[DP)0GKAKIE)P=O29THU6NF
AO^J/.FT-8>1V0B00=F=#.)7I[RT)PXe^-^[^E3YF/B\+)_;Z9IbYZI@67<;#]@A
]c6HC-+3C=]V#>14P4aI3cVJe<H;9Q_/4/MR@S1VTYCW&T[3fH#P)9W;BPP]IL>a
c>gY+_e963^);FQ\^\WF.-OKZ)TeRZaI78QcMaA0c>>>c,NW[S_FbeEL=?e1+e23
4ZYKcJ&V_PaJNH@]J)3GXcZF/#6[+\(c6b3@(f-1OCW&?V2B.fWS<eZ[ZU/4f#<Z
WTMBA>,Gg4#YcDfdV9))U^g7:]d3R0D8]L+;8,[RHc58Q7fgSS=.<#(8YD:50GeX
\2,.AD^_bMYHU?RW,C6\ZYY+0O<fAF:KV3BI#^TCF,A_?JC)Q#&_[,-S5[QKEfY1
YRWL?S7U6aUgW+a=]_RcRI\U8/6MV14C+&C.CVSP(FBQb/0.>?E)C3WPOLM,V/?3
=F);<LbP7TNN>>M[@^;:aEUT#b--+-O7Hb:1?5eV#:J6R\3>MH;(?dS0A?/D,@F,
=d6A<5QeX&E=ad>S.=AU;XO^>TRA,]VUP.Qg=g/aE(P=Lcc<DA3:#Rb>N,e9NcUJ
bN7F+g<D,HM64B[MbJ]:77R)2XK7a_4-YOM)KXgXN^=(L/3A#]>VN(EA[-f.d<)8
M5)^eVW.)SL72V^GTTc_CLHD\IYO&4^QX7Mb5g@4d9OD#WR)5;B>COa0>Ed?XB(b
<PUMPFAZB+F6<\&Z\dE/YRS2#Q\+JB-H&)e>&d+6_&.gNOO^)U+>V5F.:=9(/H>G
IaA:G:+H8NA&)bZU31+Og,_ZK(_81.a6C&Wd2AM>a</:PLD.VZd[bK\-J+df5[LW
]BD?ZBCbW+GePG0T>C-fOXO5(#Me352N3?9-eb:EF<>@-#&1=G5QDNRZ+.-d=6L4
/@567UB.=&e#c&&(#?cK_89f/P?\]XU567P9P^T54.PKO6I26;V&1e&<Y>1\3(^^
fNe>eE3gQgU1+D;_]_c?QL#Y?FH4@<_\G.+H61S^XY=#WE5fYMb_6\C6?S[S6:D?
6OGfPCd:-DgJ)8a>UUSK<L>_W,Ae\Me;]73f@b?6c_c-.V_SUEJ;4^E/20>Ge=U;
\37?e+^+0)DURDX](=ZHT:RfS/@>?O/(d>,1VD_R,\ddPS1^0VJ9+A(OP/\LSa2[
;3NG7;QL(U9g71V6H&+&_(G__3]NCGH^,H02HA:XPO.<Ic<O=R1I#XPBGR-R2a3_
f=e3NaW2&_fCB9/S_agKc,T@C?APUCK(,LTGK+N8U;,IXcFC<YU.bXDP5@Tb<e)]
8;PXXfQ(UZ52=&:KMS;7<&_P]cW:Z\+PRKI]KC^RRD65T5E7]N+B9F7]Gf,6LXS:
]O706#J^@\E64IP[IFZ3[[+W<B@@AP\]&_21-UG;W_(UbW):>A_Wg?O[cW60#P9C
>O#a#+_O/ae3d:/W3:2C+IN+RgaBRb,0?121\;Jc??@YgPMbg^X?AEQ4g=VVeBNA
C4B<cEedWIP4c\8F<:X&gfS?77Y5[Qf,d8<?TK.SP<g85]VW5:M3E?MG((I\]N3a
9J^?(B1SQK5X2;-Y=[+]XU/GfA(A(-f2,I^B70e++EP:7VN@LL6H/9KL\&#_Cac_
9FK2\KQQ\0^?g2dWV1+<_JI4:8Z@6Hfb3SJNaOB9HWF+;ZUQ-)\eC[MA2Y#V/e]2
EIcLe7<S).Y<SKR5bIf#N^f4BdTMUN)\3)\aY^?=0Y48F.^1.DPfNO3>Z+LRF\CH
=]J90;LZVPA#N9WIaS>d\45MM-WcV[6fS_;b/OfKVI=<X=J^@H5DS(I5dQbZR\=Y
X__-L4L8RQ[&g0]KP1\f(HQXb[6=+F.W>.I,4e]#@@aKG_G<Q)KW8ZN)IdOEC&K9
P,6\Q4_L]]NR[)HY\U)M_4?#AeCT7e:JF=<NW0?ZTEP/&:f,#d@84e5M7?fDc#76
fMIX/g<FYU<O.]YF==\<7^H>@:R#,0O^AC27=d3b&UA\:,?\0,5LQK^S5W,-/J5R
c[7K#GKB+4RR>dO0AVUC3MTb\?E17K_DId@0cJA<ZGNc]J)4Y@.fH&b8;JU?;&&+
Wg0A<6D4Wb4/Sfbc@2SRb>IT,UX1Uf3LA_]Fg?4a46G9O\F505&Ia.D1)^2af9)U
aE7Z5IWO/]TA#D#eWL)&NL-WUe75BQP:JJ?V:YBg@IL;PCL4cR9eW:#K3PVX:TVJ
_VP919ZJNUH.5:Y#+b<>60<]WL&AG8S(S3P,TM3S_.bD_TFK0G<\7&8Y]KgGHPO+
J&ZHgeO7U1;dPgdH8VTNb>S2C5B,NN15^U>=8.KUT^3?+/SX/MBV:NIQcTdRC)#M
R6,?\@QPUM6L<RK(,<)g4X\ZCa77^]XfaF<9+N[^;QR@D0:2IM4O.#SQ80KXMIZH
=[LcV3<PbE.1Vb?4(3>;ed[[RXVNPL.<8;-fa?8f4)/8Ya4&9:N<EEZ#^B]Fbc6)
7@F=@>5BP;/4-gXTJGcAOAcfd-3?;.[L)5FB,0>C3ag<@8QHA<5#(U>;[U-8+L_#
RS>ZLL^:-J8dSX&5K<8S_,3)C-3\AVS\/=6eEIfPd?&Z9]=,1H(^\;T2]5.+6KBN
04<dP40\B#8X7J6N\-FW(G&CV&73F\+FZJfc1C=_5N?_NZSQ<Z?=O#6,EK/KZ:6[
/bPV0ee;L54\0Y0b:0[BUCbUF\#=M546:c#.A-B\N2TFd8fge\CP-^e7J<K:ZD@&
U2?d1dLgL)M5^1W^b:GY60;O?M+C\N[LaJf<F,H\Q8,&.a(D<//DT6:Q-+[386/S
M,MSLOC]==Xc8MF\NdBZfJQ>EI)M6G/J42BV+eTNR5_)Y&OQOX#CCAP[DVYUU.?N
X:?5T@8=bO;+3GKN?7b3.UG;a]Q9.OH44I#@[MR6X;@BUDXIA=[3@8>E8I8S\)de
a7L1]Z+6CT=aSG.a:g=JHCGH;EG2V](4gXN7WM3A5W=e8103#\?I:[,5:5+)e\Sc
c[gKZ=/.,)<U-Q4&7\,I6HKI:H32gQ-3&?>d[9I^7QZ_@ET6#2Y4/f,?WOZg[fb2
K\Cb+&K/cbEZ_HBDW[?6Hf+Y.L:aBCDSCXgZg0g_O,PSa\E;/;:DT-^a+S4C(C\f
2+X+dQ_^O2;,=-X#UX5L_MN<UO2?:DB4T+N#c<b(SL99[5WeRH:]_27@N,61dWO;
EO2P9<IGQ+4Ed@g(KSJIH>Jc\JO7;#)c1Ib&9.)K&2<^&c;<2E_bB[=)bL+Z(.6\
+>YB<.8A&[#A,G=]7LKRaP0I]3?-XM.+(M[bX)9:04G.eI=\YWE?aY7PXP<G=]J(
6<&3f1./Mg/=C(F(J5a34X2e0IU^6ZZC4:6d5bJ8T&6Y^SQ&0/df89\]+&\#Y=Y_
?(24@cV_/Z#=4Y\?D>+6gaeJ3)GZLEPQ^+0MZO)8;1?#3L)U6^Le)1TE+O?cF8e7
)=&QA>gM)CUG]fAZ#&#=[U3\#P5EZbXK).BWRF5?19/\BL^9,BK_(bI,<2LaP5Xb
\,)AUHe]K[@P,.]J()X;B[^a/TOX(.+JB)/De2XYV(Oe]FQE,O;LF]LSBKdI(<_-
Z^_0BP.6[D8PE1W_YS/S=:cGb=Od.IXXD-2UG\/-\A2<f2)0c22TP#@cTNa3V#OG
_+T37R<25cW:2@<eA.4Uc8[OKMB;41gS4)cd3L1WFMaK>((,c3TS@^dE<,_E=c4H
Q[e;?#&<EFJBLS2dCGB=81<cAb5N(A^ZXQ:a1TDbJJ:E)A)KS)D<^f[+4?M1<[I^
<QXQXASJ&fPJZEg1@+d\UB6,3fg>;[B.?JfOQ]_+HE5[_H,4HScS<150#OUWc7>=
gAAC..b9bDU(4Ie+DWU>=W0_N\IY)aU[BZd/49PLYFR1U,N4De/S,^CWF./O0\4d
P;AF-<#)5MD&EMa9:<<<1bY-]<5Q1eTW=WcEPbQg7Y0PgP7/4YG.BP^).MW&gbY/
4Z=P&a/f<a^\14Y:=U-RY9.VBZNCg+;3cNT/dN)c;C8IYB<UUE5[A_8XI6=BI7JE
Z8&McTPG89)A08c+2W_B;&f1[><2GO981cYW9@,4LC+8cTe8_&U2H8G4BfS4D&<-
5=P1##K<C)8EXEbDF7Z)0K4V=^a;-dWY>8;&<eMb_\N+g/?RLAXNH=\f??@gdW-6
](+X0T=V_@e=,&Y=_F#8T5SQdUMZ^DCW?T05eB,aG=5>:RTHPZ16(EeEN4C7d>-3
fM;V+X48[gI6)J3D?gOF4+B#H^9ITbZ6Ab+NRB-SUUVP.B-:FdX9bVDL5OdeZ0K5
2ef0.IV0\9BV7d,(Q-T9ORJ3XOL0[<QRHOC/N97B.[&W^OgM((+gcRISaI>EDX4(
&NFI>G5E:-[M^OLNGe@^1[C7U7+&d&PHV)+/A]]Z_1^>AY][Y,,=XL@0(_d1/2=Y
QJ@_-86HA/:U2L<0W^=>^SY4MNNgdDZMGTG],2YUX:-OGJ[73b,O(&@0I$
`endprotected
endmodule
